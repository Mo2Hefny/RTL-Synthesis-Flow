module floating_point_alu (overflow,
    sel,
    a,
    b,
    result);
 output overflow;
 input sel;
 input [31:0] a;
 input [31:0] b;
 output [31:0] result;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;

 sky130_fd_sc_hd__inv_12 _05350_ (.A(net65),
    .Y(_05339_));
 sky130_fd_sc_hd__inv_6 _05351_ (.A(net16),
    .Y(_00000_));
 sky130_fd_sc_hd__clkinv_4 _05352_ (.A(net19),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_6 _05353_ (.A(net12),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_8 _05354_ (.A(net1),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_6 _05355_ (.A(net26),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_6 _05356_ (.A(net23),
    .Y(_00055_));
 sky130_fd_sc_hd__clkinv_8 _05357_ (.A(net28),
    .Y(_00066_));
 sky130_fd_sc_hd__clkinv_8 _05358_ (.A(net27),
    .Y(_00077_));
 sky130_fd_sc_hd__inv_6 _05359_ (.A(net30),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_6 _05360_ (.A(net29),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_8 _05361_ (.A(net32),
    .Y(_00110_));
 sky130_fd_sc_hd__clkinv_8 _05362_ (.A(net31),
    .Y(_00121_));
 sky130_fd_sc_hd__inv_8 _05363_ (.A(net3),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_8 _05364_ (.A(net2),
    .Y(_00143_));
 sky130_fd_sc_hd__clkinv_8 _05365_ (.A(net5),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_8 _05366_ (.A(net4),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_8 _05367_ (.A(net7),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_8 _05368_ (.A(net6),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_6 _05369_ (.A(net9),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_8 _05370_ (.A(net8),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_6 _05371_ (.A(net11),
    .Y(_00220_));
 sky130_fd_sc_hd__clkinv_8 _05372_ (.A(net10),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_6 _05373_ (.A(net14),
    .Y(_00242_));
 sky130_fd_sc_hd__clkinv_8 _05374_ (.A(net13),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_8 _05375_ (.A(net15),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _05376_ (.A(net50),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _05377_ (.A(net53),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _05378_ (.A(net56),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _05379_ (.A(net44),
    .Y(_00308_));
 sky130_fd_sc_hd__inv_2 _05380_ (.A(net33),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _05381_ (.A(net58),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_16 _05382_ (.A(net55),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_16 _05383_ (.A(net60),
    .Y(_00352_));
 sky130_fd_sc_hd__clkinv_4 _05384_ (.A(net59),
    .Y(_00363_));
 sky130_fd_sc_hd__clkinv_8 _05385_ (.A(net62),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_6 _05386_ (.A(net61),
    .Y(_00385_));
 sky130_fd_sc_hd__clkinv_16 _05387_ (.A(net63),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_16 _05388_ (.A(net35),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_2 _05389_ (.A(net34),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_4 _05390_ (.A(net36),
    .Y(_00429_));
 sky130_fd_sc_hd__clkinv_8 _05391_ (.A(net39),
    .Y(_00440_));
 sky130_fd_sc_hd__inv_16 _05392_ (.A(net41),
    .Y(_00451_));
 sky130_fd_sc_hd__inv_8 _05393_ (.A(net43),
    .Y(_00462_));
 sky130_fd_sc_hd__clkinv_8 _05394_ (.A(net42),
    .Y(_00473_));
 sky130_fd_sc_hd__clkinv_8 _05395_ (.A(net46),
    .Y(_00484_));
 sky130_fd_sc_hd__and4_1 _05396_ (.A(net53),
    .B(net52),
    .C(net54),
    .D(net56),
    .X(_00495_));
 sky130_fd_sc_hd__and3_1 _05397_ (.A(net49),
    .B(net48),
    .C(net51),
    .X(_00506_));
 sky130_fd_sc_hd__and3_2 _05398_ (.A(net50),
    .B(_00495_),
    .C(_00506_),
    .X(_00517_));
 sky130_fd_sc_hd__or4_1 _05399_ (.A(net41),
    .B(net42),
    .C(net46),
    .D(net47),
    .X(_00528_));
 sky130_fd_sc_hd__nor4_1 _05400_ (.A(net40),
    .B(net43),
    .C(net45),
    .D(_00528_),
    .Y(_00539_));
 sky130_fd_sc_hd__and4b_1 _05401_ (.A_N(net64),
    .B(_00396_),
    .C(_00407_),
    .D(_00418_),
    .X(_00550_));
 sky130_fd_sc_hd__nor4_1 _05402_ (.A(net37),
    .B(net36),
    .C(net39),
    .D(net38),
    .Y(_00561_));
 sky130_fd_sc_hd__and3_2 _05403_ (.A(_00539_),
    .B(_00550_),
    .C(_00561_),
    .X(_00572_));
 sky130_fd_sc_hd__and4_2 _05404_ (.A(_00308_),
    .B(_00319_),
    .C(_00330_),
    .D(_00341_),
    .X(_00583_));
 sky130_fd_sc_hd__and4_2 _05405_ (.A(_00352_),
    .B(_00363_),
    .C(_00374_),
    .D(_00385_),
    .X(_00594_));
 sky130_fd_sc_hd__nand3_1 _05406_ (.A(_00572_),
    .B(_00583_),
    .C(_00594_),
    .Y(_00605_));
 sky130_fd_sc_hd__and4_1 _05407_ (.A(net21),
    .B(net20),
    .C(net22),
    .D(net24),
    .X(_00616_));
 sky130_fd_sc_hd__and3_1 _05408_ (.A(net17),
    .B(net16),
    .C(net19),
    .X(_00627_));
 sky130_fd_sc_hd__and3_2 _05409_ (.A(net18),
    .B(_00616_),
    .C(_00627_),
    .X(_00638_));
 sky130_fd_sc_hd__or4_1 _05410_ (.A(net9),
    .B(net10),
    .C(net14),
    .D(net15),
    .X(_00649_));
 sky130_fd_sc_hd__and4b_1 _05411_ (.A_N(_00649_),
    .B(_00253_),
    .C(_00220_),
    .D(_00209_),
    .X(_00660_));
 sky130_fd_sc_hd__and4_1 _05412_ (.A(_00110_),
    .B(_00121_),
    .C(_00132_),
    .D(_00143_),
    .X(_00671_));
 sky130_fd_sc_hd__and4_1 _05413_ (.A(_00154_),
    .B(_00165_),
    .C(_00176_),
    .D(_00187_),
    .X(_00682_));
 sky130_fd_sc_hd__and3_1 _05414_ (.A(_00660_),
    .B(_00671_),
    .C(_00682_),
    .X(_00693_));
 sky130_fd_sc_hd__and4_1 _05415_ (.A(_00022_),
    .B(_00033_),
    .C(_00044_),
    .D(_00055_),
    .X(_00704_));
 sky130_fd_sc_hd__and4_1 _05416_ (.A(_00066_),
    .B(_00077_),
    .C(_00088_),
    .D(_00099_),
    .X(_00715_));
 sky130_fd_sc_hd__nand3_4 _05417_ (.A(_00693_),
    .B(_00704_),
    .C(_00715_),
    .Y(_00726_));
 sky130_fd_sc_hd__inv_2 _05418_ (.A(_00726_),
    .Y(_00737_));
 sky130_fd_sc_hd__a22oi_2 _05419_ (.A1(_00517_),
    .A2(_00605_),
    .B1(_00726_),
    .B2(_00638_),
    .Y(_00748_));
 sky130_fd_sc_hd__nor3_1 _05420_ (.A(net53),
    .B(net52),
    .C(net54),
    .Y(_00759_));
 sky130_fd_sc_hd__nor3_2 _05421_ (.A(net49),
    .B(net48),
    .C(net51),
    .Y(_00770_));
 sky130_fd_sc_hd__and4_4 _05422_ (.A(_00759_),
    .B(_00770_),
    .C(_00275_),
    .D(_00297_),
    .X(_00781_));
 sky130_fd_sc_hd__nand4_4 _05423_ (.A(_00759_),
    .B(_00770_),
    .C(_00275_),
    .D(_00297_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand2_2 _05424_ (.A(_00638_),
    .B(_00737_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_1 _05425_ (.A(net20),
    .B(net22),
    .Y(_00814_));
 sky130_fd_sc_hd__nor2_1 _05426_ (.A(net21),
    .B(net24),
    .Y(_00825_));
 sky130_fd_sc_hd__nor4_4 _05427_ (.A(net21),
    .B(net20),
    .C(net22),
    .D(net24),
    .Y(_00836_));
 sky130_fd_sc_hd__nor3_4 _05428_ (.A(net17),
    .B(net19),
    .C(net18),
    .Y(_00847_));
 sky130_fd_sc_hd__nor4_4 _05429_ (.A(net17),
    .B(net16),
    .C(net19),
    .D(net18),
    .Y(_00858_));
 sky130_fd_sc_hd__and3_4 _05430_ (.A(net118),
    .B(_00847_),
    .C(_00000_),
    .X(_00869_));
 sky130_fd_sc_hd__nand4_4 _05431_ (.A(_00814_),
    .B(_00825_),
    .C(_00847_),
    .D(_00000_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand4_2 _05432_ (.A(_00517_),
    .B(_00572_),
    .C(_00583_),
    .D(_00594_),
    .Y(_00891_));
 sky130_fd_sc_hd__or3_1 _05433_ (.A(_00726_),
    .B(_00880_),
    .C(_00891_),
    .X(_00902_));
 sky130_fd_sc_hd__o31a_1 _05434_ (.A1(_00605_),
    .A2(_00792_),
    .A3(_00803_),
    .B1(_00902_),
    .X(_00913_));
 sky130_fd_sc_hd__nand2_1 _05435_ (.A(_00748_),
    .B(_00913_),
    .Y(_00924_));
 sky130_fd_sc_hd__or2_1 _05436_ (.A(_05339_),
    .B(_00924_),
    .X(_00935_));
 sky130_fd_sc_hd__nor2_8 _05437_ (.A(net16),
    .B(net48),
    .Y(_00946_));
 sky130_fd_sc_hd__or2_4 _05438_ (.A(net16),
    .B(net48),
    .X(_00957_));
 sky130_fd_sc_hd__and2b_1 _05439_ (.A_N(net17),
    .B(net49),
    .X(_00968_));
 sky130_fd_sc_hd__nand2b_1 _05440_ (.A_N(net17),
    .B(net49),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2b_2 _05441_ (.A_N(net49),
    .B(net17),
    .Y(_00990_));
 sky130_fd_sc_hd__nand2_4 _05442_ (.A(_00979_),
    .B(_00990_),
    .Y(_01001_));
 sky130_fd_sc_hd__xnor2_4 _05443_ (.A(net17),
    .B(net49),
    .Y(_01012_));
 sky130_fd_sc_hd__nor2_4 _05444_ (.A(net18),
    .B(_00275_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2b_1 _05445_ (.A_N(net18),
    .B(net50),
    .Y(_01034_));
 sky130_fd_sc_hd__and2_1 _05446_ (.A(_00275_),
    .B(net18),
    .X(_01045_));
 sky130_fd_sc_hd__nand2b_2 _05447_ (.A_N(net50),
    .B(net18),
    .Y(_01056_));
 sky130_fd_sc_hd__nand2_1 _05448_ (.A(_01034_),
    .B(_01056_),
    .Y(_01067_));
 sky130_fd_sc_hd__o211ai_1 _05449_ (.A1(_01023_),
    .A2(_01045_),
    .B1(net17),
    .C1(net49),
    .Y(_01078_));
 sky130_fd_sc_hd__a211o_1 _05450_ (.A1(net17),
    .A2(net49),
    .B1(_01023_),
    .C1(_01045_),
    .X(_01089_));
 sky130_fd_sc_hd__o221a_1 _05451_ (.A1(net16),
    .A2(net48),
    .B1(_01023_),
    .B2(_01045_),
    .C1(_01001_),
    .X(_01100_));
 sky130_fd_sc_hd__nand2_1 _05452_ (.A(_00011_),
    .B(net51),
    .Y(_01111_));
 sky130_fd_sc_hd__or2_2 _05453_ (.A(net51),
    .B(_00011_),
    .X(_01122_));
 sky130_fd_sc_hd__xnor2_4 _05454_ (.A(net19),
    .B(net51),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_2 _05455_ (.A(_01111_),
    .B(_01122_),
    .Y(_01144_));
 sky130_fd_sc_hd__or3b_1 _05456_ (.A(_01133_),
    .B(_00275_),
    .C_N(net18),
    .X(_01155_));
 sky130_fd_sc_hd__a21o_1 _05457_ (.A1(net18),
    .A2(net50),
    .B1(_01144_),
    .X(_01166_));
 sky130_fd_sc_hd__nand2_1 _05458_ (.A(_01155_),
    .B(_01166_),
    .Y(_01177_));
 sky130_fd_sc_hd__a31o_2 _05459_ (.A1(net17),
    .A2(net49),
    .A3(_01067_),
    .B1(_01100_),
    .X(_01188_));
 sky130_fd_sc_hd__a21boi_2 _05460_ (.A1(_01166_),
    .A2(_01188_),
    .B1_N(_01155_),
    .Y(_01199_));
 sky130_fd_sc_hd__and2_1 _05461_ (.A(net20),
    .B(net52),
    .X(_01210_));
 sky130_fd_sc_hd__nor2_1 _05462_ (.A(net20),
    .B(net52),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_2 _05463_ (.A(_01210_),
    .B(_01221_),
    .Y(_01232_));
 sky130_fd_sc_hd__or2_1 _05464_ (.A(_01210_),
    .B(_01221_),
    .X(_01243_));
 sky130_fd_sc_hd__and3_1 _05465_ (.A(net19),
    .B(net51),
    .C(_01232_),
    .X(_01254_));
 sky130_fd_sc_hd__o2bb2a_1 _05466_ (.A1_N(net19),
    .A2_N(net51),
    .B1(_01210_),
    .B2(_01221_),
    .X(_01265_));
 sky130_fd_sc_hd__or2_1 _05467_ (.A(_01254_),
    .B(_01265_),
    .X(_01276_));
 sky130_fd_sc_hd__and2_1 _05468_ (.A(net21),
    .B(net53),
    .X(_01287_));
 sky130_fd_sc_hd__nand2_4 _05469_ (.A(net21),
    .B(net53),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_2 _05470_ (.A(net21),
    .B(net53),
    .Y(_01309_));
 sky130_fd_sc_hd__or2_4 _05471_ (.A(net21),
    .B(net53),
    .X(_01320_));
 sky130_fd_sc_hd__o2bb2a_1 _05472_ (.A1_N(net20),
    .A2_N(net52),
    .B1(_01287_),
    .B2(_01309_),
    .X(_01331_));
 sky130_fd_sc_hd__and3_1 _05473_ (.A(_01320_),
    .B(_01210_),
    .C(_01298_),
    .X(_01342_));
 sky130_fd_sc_hd__or2_1 _05474_ (.A(_01331_),
    .B(_01342_),
    .X(_01353_));
 sky130_fd_sc_hd__or4_4 _05475_ (.A(_01254_),
    .B(_01265_),
    .C(_01331_),
    .D(_01342_),
    .X(_01364_));
 sky130_fd_sc_hd__inv_2 _05476_ (.A(_01364_),
    .Y(_01375_));
 sky130_fd_sc_hd__a31o_1 _05477_ (.A1(_01254_),
    .A2(_01298_),
    .A3(_01320_),
    .B1(_01342_),
    .X(_01386_));
 sky130_fd_sc_hd__o21ba_1 _05478_ (.A1(_01199_),
    .A2(_01364_),
    .B1_N(_01386_),
    .X(_01397_));
 sky130_fd_sc_hd__and2b_1 _05479_ (.A_N(net22),
    .B(net54),
    .X(_01408_));
 sky130_fd_sc_hd__nand2b_2 _05480_ (.A_N(net22),
    .B(net54),
    .Y(_01419_));
 sky130_fd_sc_hd__and2b_2 _05481_ (.A_N(net54),
    .B(net22),
    .X(_01430_));
 sky130_fd_sc_hd__nand2b_2 _05482_ (.A_N(net54),
    .B(net22),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _05483_ (.A(_01408_),
    .B(_01430_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_4 _05484_ (.A(_01419_),
    .B(_01441_),
    .Y(_01463_));
 sky130_fd_sc_hd__xor2_1 _05485_ (.A(_01298_),
    .B(_01463_),
    .X(_01474_));
 sky130_fd_sc_hd__nor2_1 _05486_ (.A(_01474_),
    .B(_01397_),
    .Y(_01485_));
 sky130_fd_sc_hd__and2_1 _05487_ (.A(_01397_),
    .B(_01474_),
    .X(_01496_));
 sky130_fd_sc_hd__nor2_1 _05488_ (.A(_01485_),
    .B(_01496_),
    .Y(_01507_));
 sky130_fd_sc_hd__inv_2 _05489_ (.A(_01507_),
    .Y(_01518_));
 sky130_fd_sc_hd__and2_4 _05490_ (.A(net16),
    .B(net48),
    .X(_01529_));
 sky130_fd_sc_hd__nand2_4 _05491_ (.A(net16),
    .B(net48),
    .Y(_01540_));
 sky130_fd_sc_hd__nor2_8 _05492_ (.A(_00946_),
    .B(_01529_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_8 _05493_ (.A(_00957_),
    .B(_01540_),
    .Y(_01562_));
 sky130_fd_sc_hd__and2_1 _05494_ (.A(net15),
    .B(net47),
    .X(_01573_));
 sky130_fd_sc_hd__nand2_1 _05495_ (.A(net15),
    .B(net47),
    .Y(_01584_));
 sky130_fd_sc_hd__a22o_1 _05496_ (.A1(_00880_),
    .A2(net47),
    .B1(net15),
    .B2(_00792_),
    .X(_01595_));
 sky130_fd_sc_hd__o31a_1 _05497_ (.A1(_01584_),
    .A2(_00869_),
    .A3(_00781_),
    .B1(_01595_),
    .X(_01606_));
 sky130_fd_sc_hd__and3_1 _05498_ (.A(_00880_),
    .B(_01573_),
    .C(net46),
    .X(_01617_));
 sky130_fd_sc_hd__o2bb2a_1 _05499_ (.A1_N(net15),
    .A2_N(net47),
    .B1(_00484_),
    .B2(_00869_),
    .X(_01628_));
 sky130_fd_sc_hd__a22o_1 _05500_ (.A1(net15),
    .A2(net47),
    .B1(_00880_),
    .B2(net46),
    .X(_01639_));
 sky130_fd_sc_hd__and4b_1 _05501_ (.A_N(_01617_),
    .B(net14),
    .C(_00792_),
    .D(_01639_),
    .X(_01650_));
 sky130_fd_sc_hd__a31o_1 _05502_ (.A1(_01639_),
    .A2(net14),
    .A3(_00792_),
    .B1(_01617_),
    .X(_01661_));
 sky130_fd_sc_hd__o311a_1 _05503_ (.A1(_00781_),
    .A2(_00869_),
    .A3(_01584_),
    .B1(_01595_),
    .C1(_01661_),
    .X(_01672_));
 sky130_fd_sc_hd__or4b_2 _05504_ (.A(_00781_),
    .B(_00869_),
    .C(_01573_),
    .D_N(_01672_),
    .X(_01683_));
 sky130_fd_sc_hd__o31a_4 _05505_ (.A1(_00781_),
    .A2(_00869_),
    .A3(_01584_),
    .B1(_01683_),
    .X(_01694_));
 sky130_fd_sc_hd__o22a_1 _05506_ (.A1(_00242_),
    .A2(_00781_),
    .B1(_01617_),
    .B2(_01628_),
    .X(_01705_));
 sky130_fd_sc_hd__and3_1 _05507_ (.A(net14),
    .B(net46),
    .C(_01573_),
    .X(_01716_));
 sky130_fd_sc_hd__a22oi_1 _05508_ (.A1(net15),
    .A2(net46),
    .B1(net47),
    .B2(net14),
    .Y(_01727_));
 sky130_fd_sc_hd__a22o_1 _05509_ (.A1(net15),
    .A2(net46),
    .B1(net47),
    .B2(net14),
    .X(_01738_));
 sky130_fd_sc_hd__and4b_1 _05510_ (.A_N(_01716_),
    .B(net13),
    .C(_00792_),
    .D(_01738_),
    .X(_01749_));
 sky130_fd_sc_hd__a31o_1 _05511_ (.A1(net13),
    .A2(_00792_),
    .A3(_01738_),
    .B1(_01716_),
    .X(_01760_));
 sky130_fd_sc_hd__nor2_1 _05512_ (.A(_00264_),
    .B(_00462_),
    .Y(_01771_));
 sky130_fd_sc_hd__o22a_1 _05513_ (.A1(_01716_),
    .A2(_01727_),
    .B1(_00253_),
    .B2(_00781_),
    .X(_01782_));
 sky130_fd_sc_hd__nor2_1 _05514_ (.A(_01749_),
    .B(_01782_),
    .Y(_01793_));
 sky130_fd_sc_hd__or3b_1 _05515_ (.A(_00869_),
    .B(_01771_),
    .C_N(net45),
    .X(_01804_));
 sky130_fd_sc_hd__o2111a_1 _05516_ (.A1(_00264_),
    .A2(_00462_),
    .B1(net45),
    .C1(_00880_),
    .D1(_01793_),
    .X(_01815_));
 sky130_fd_sc_hd__o2111a_1 _05517_ (.A1(_01771_),
    .A2(_01793_),
    .B1(net45),
    .C1(_00880_),
    .D1(_01760_),
    .X(_01826_));
 sky130_fd_sc_hd__a311o_1 _05518_ (.A1(net45),
    .A2(_00880_),
    .A3(_01771_),
    .B1(_01760_),
    .C1(_01815_),
    .X(_01837_));
 sky130_fd_sc_hd__nand2b_1 _05519_ (.A_N(_01826_),
    .B(_01837_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor3_1 _05520_ (.A(_01650_),
    .B(_01705_),
    .C(_01848_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _05521_ (.A(_01606_),
    .B(_01661_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _05522_ (.A(_01672_),
    .B(_01870_),
    .Y(_01881_));
 sky130_fd_sc_hd__or4b_1 _05523_ (.A(_01650_),
    .B(_01705_),
    .C(_01848_),
    .D_N(_01881_),
    .X(_01892_));
 sky130_fd_sc_hd__or2_1 _05524_ (.A(_01859_),
    .B(_01881_),
    .X(_01903_));
 sky130_fd_sc_hd__o21ai_2 _05525_ (.A1(_01826_),
    .A2(_01859_),
    .B1(_01881_),
    .Y(_01914_));
 sky130_fd_sc_hd__inv_2 _05526_ (.A(_01914_),
    .Y(_01925_));
 sky130_fd_sc_hd__a31o_1 _05527_ (.A1(_00792_),
    .A2(_00880_),
    .A3(_01584_),
    .B1(_01672_),
    .X(_01936_));
 sky130_fd_sc_hd__nand2_2 _05528_ (.A(_01683_),
    .B(_01936_),
    .Y(_01947_));
 sky130_fd_sc_hd__or2_4 _05529_ (.A(_01947_),
    .B(_01914_),
    .X(_01958_));
 sky130_fd_sc_hd__xor2_1 _05530_ (.A(_01793_),
    .B(_01804_),
    .X(_01969_));
 sky130_fd_sc_hd__and4_1 _05531_ (.A(net14),
    .B(net13),
    .C(net46),
    .D(net47),
    .X(_01980_));
 sky130_fd_sc_hd__a22oi_1 _05532_ (.A1(net14),
    .A2(net46),
    .B1(net47),
    .B2(net13),
    .Y(_01991_));
 sky130_fd_sc_hd__a22o_1 _05533_ (.A1(net14),
    .A2(net46),
    .B1(net47),
    .B2(net13),
    .X(_02002_));
 sky130_fd_sc_hd__a31o_1 _05534_ (.A1(_00792_),
    .A2(_02002_),
    .A3(net11),
    .B1(_01980_),
    .X(_02013_));
 sky130_fd_sc_hd__a211oi_1 _05535_ (.A1(_00792_),
    .A2(net11),
    .B1(_01991_),
    .C1(_01980_),
    .Y(_02024_));
 sky130_fd_sc_hd__o211a_1 _05536_ (.A1(_01980_),
    .A2(_01991_),
    .B1(net11),
    .C1(_00792_),
    .X(_02035_));
 sky130_fd_sc_hd__nor2_1 _05537_ (.A(_02024_),
    .B(_02035_),
    .Y(_02046_));
 sky130_fd_sc_hd__o2bb2a_1 _05538_ (.A1_N(net15),
    .A2_N(net45),
    .B1(_00462_),
    .B2(_00869_),
    .X(_02057_));
 sky130_fd_sc_hd__a31oi_1 _05539_ (.A1(net45),
    .A2(_00880_),
    .A3(_01771_),
    .B1(_02057_),
    .Y(_02068_));
 sky130_fd_sc_hd__and4_1 _05540_ (.A(_00880_),
    .B(net42),
    .C(net43),
    .D(net15),
    .X(_02079_));
 sky130_fd_sc_hd__o22a_1 _05541_ (.A1(_00264_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00869_),
    .X(_02090_));
 sky130_fd_sc_hd__and4bb_1 _05542_ (.A_N(_02079_),
    .B_N(_02090_),
    .C(net14),
    .D(net45),
    .X(_02101_));
 sky130_fd_sc_hd__o21a_1 _05543_ (.A1(_02079_),
    .A2(_02101_),
    .B1(_02068_),
    .X(_02112_));
 sky130_fd_sc_hd__or3_1 _05544_ (.A(_02068_),
    .B(_02079_),
    .C(_02101_),
    .X(_02123_));
 sky130_fd_sc_hd__nand2b_1 _05545_ (.A_N(_02112_),
    .B(_02123_),
    .Y(_02134_));
 sky130_fd_sc_hd__xnor2_1 _05546_ (.A(_02046_),
    .B(_02134_),
    .Y(_02145_));
 sky130_fd_sc_hd__and2_1 _05547_ (.A(net15),
    .B(net40),
    .X(_02156_));
 sky130_fd_sc_hd__and3_1 _05548_ (.A(_00880_),
    .B(_02156_),
    .C(net41),
    .X(_02167_));
 sky130_fd_sc_hd__and3_1 _05549_ (.A(net14),
    .B(net42),
    .C(_01771_),
    .X(_02178_));
 sky130_fd_sc_hd__o22a_1 _05550_ (.A1(_00242_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00264_),
    .X(_02189_));
 sky130_fd_sc_hd__and4bb_1 _05551_ (.A_N(_02178_),
    .B_N(_02189_),
    .C(net13),
    .D(net45),
    .X(_02200_));
 sky130_fd_sc_hd__o2bb2a_1 _05552_ (.A1_N(net14),
    .A2_N(net45),
    .B1(_02079_),
    .B2(_02090_),
    .X(_02211_));
 sky130_fd_sc_hd__or2_1 _05553_ (.A(_02101_),
    .B(_02211_),
    .X(_02222_));
 sky130_fd_sc_hd__o21bai_1 _05554_ (.A1(_02178_),
    .A2(_02200_),
    .B1_N(_02222_),
    .Y(_02233_));
 sky130_fd_sc_hd__or3b_1 _05555_ (.A(_02178_),
    .B(_02200_),
    .C_N(_02222_),
    .X(_02244_));
 sky130_fd_sc_hd__nand2_1 _05556_ (.A(_02233_),
    .B(_02244_),
    .Y(_02255_));
 sky130_fd_sc_hd__a22oi_1 _05557_ (.A1(net13),
    .A2(net46),
    .B1(net47),
    .B2(net11),
    .Y(_02266_));
 sky130_fd_sc_hd__and4_1 _05558_ (.A(net11),
    .B(net13),
    .C(net46),
    .D(net47),
    .X(_02277_));
 sky130_fd_sc_hd__or4_1 _05559_ (.A(_02266_),
    .B(_00231_),
    .C(_00781_),
    .D(_02277_),
    .X(_02288_));
 sky130_fd_sc_hd__a2bb2o_1 _05560_ (.A1_N(_02266_),
    .A2_N(_02277_),
    .B1(net10),
    .B2(net117),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_1 _05561_ (.A(_02288_),
    .B(_02299_),
    .Y(_02310_));
 sky130_fd_sc_hd__or2_1 _05562_ (.A(_02255_),
    .B(_02310_),
    .X(_02321_));
 sky130_fd_sc_hd__nand2_1 _05563_ (.A(_02255_),
    .B(_02310_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand2_1 _05564_ (.A(_02321_),
    .B(_02332_),
    .Y(_02343_));
 sky130_fd_sc_hd__or4b_2 _05565_ (.A(_00451_),
    .B(_02343_),
    .C(_00869_),
    .D_N(_02156_),
    .X(_02354_));
 sky130_fd_sc_hd__o31ai_1 _05566_ (.A1(_02024_),
    .A2(_02035_),
    .A3(_02112_),
    .B1(_02123_),
    .Y(_02365_));
 sky130_fd_sc_hd__or3_1 _05567_ (.A(_02145_),
    .B(_02354_),
    .C(_02365_),
    .X(_02376_));
 sky130_fd_sc_hd__o21ai_1 _05568_ (.A1(_02145_),
    .A2(_02354_),
    .B1(_02365_),
    .Y(_02387_));
 sky130_fd_sc_hd__and2_1 _05569_ (.A(_02376_),
    .B(_02387_),
    .X(_02398_));
 sky130_fd_sc_hd__xnor2_1 _05570_ (.A(_02013_),
    .B(_02398_),
    .Y(_02409_));
 sky130_fd_sc_hd__or2_1 _05571_ (.A(_01969_),
    .B(_02409_),
    .X(_02420_));
 sky130_fd_sc_hd__o21a_1 _05572_ (.A1(_01650_),
    .A2(_01705_),
    .B1(_01848_),
    .X(_02431_));
 sky130_fd_sc_hd__or2_1 _05573_ (.A(_01859_),
    .B(_02431_),
    .X(_02442_));
 sky130_fd_sc_hd__a21bo_1 _05574_ (.A1(_02013_),
    .A2(_02387_),
    .B1_N(_02376_),
    .X(_02453_));
 sky130_fd_sc_hd__xnor2_1 _05575_ (.A(_02420_),
    .B(_02442_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2b_1 _05576_ (.A_N(_02464_),
    .B(_02453_),
    .Y(_02475_));
 sky130_fd_sc_hd__o21ai_1 _05577_ (.A1(_02420_),
    .A2(_02442_),
    .B1(_02475_),
    .Y(_02486_));
 sky130_fd_sc_hd__a21oi_1 _05578_ (.A1(_01892_),
    .A2(_01903_),
    .B1(_01826_),
    .Y(_02497_));
 sky130_fd_sc_hd__a21oi_1 _05579_ (.A1(_01826_),
    .A2(_01881_),
    .B1(_02497_),
    .Y(_02508_));
 sky130_fd_sc_hd__nand2_1 _05580_ (.A(_02486_),
    .B(_02508_),
    .Y(_02519_));
 sky130_fd_sc_hd__inv_2 _05581_ (.A(_02519_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _05582_ (.A(_02508_),
    .B(_02486_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _05583_ (.A(_02530_),
    .B(_02541_),
    .Y(_02552_));
 sky130_fd_sc_hd__nand2b_1 _05584_ (.A_N(_02453_),
    .B(_02464_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _05585_ (.A(_02475_),
    .B(_02563_),
    .Y(_02574_));
 sky130_fd_sc_hd__nand2_1 _05586_ (.A(_01969_),
    .B(_02409_),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _05587_ (.A(_02420_),
    .B(_02585_),
    .Y(_02596_));
 sky130_fd_sc_hd__xnor2_1 _05588_ (.A(_02145_),
    .B(_02354_),
    .Y(_02607_));
 sky130_fd_sc_hd__and2b_1 _05589_ (.A_N(_02277_),
    .B(_02288_),
    .X(_02618_));
 sky130_fd_sc_hd__o2bb2a_1 _05590_ (.A1_N(net40),
    .A2_N(_00880_),
    .B1(_00264_),
    .B2(_00451_),
    .X(_02629_));
 sky130_fd_sc_hd__nor2_1 _05591_ (.A(_02167_),
    .B(_02629_),
    .Y(_02640_));
 sky130_fd_sc_hd__and3_1 _05592_ (.A(_00880_),
    .B(_02156_),
    .C(net39),
    .X(_02651_));
 sky130_fd_sc_hd__o2bb2a_1 _05593_ (.A1_N(net15),
    .A2_N(net40),
    .B1(_00440_),
    .B2(_00869_),
    .X(_02662_));
 sky130_fd_sc_hd__nor4_1 _05594_ (.A(_00242_),
    .B(_00451_),
    .C(_02651_),
    .D(_02662_),
    .Y(_02673_));
 sky130_fd_sc_hd__o21ai_2 _05595_ (.A1(_02651_),
    .A2(_02673_),
    .B1(_02640_),
    .Y(_02684_));
 sky130_fd_sc_hd__a2111oi_1 _05596_ (.A1(net15),
    .A2(net40),
    .B1(_00869_),
    .C1(_02684_),
    .D1(_00451_),
    .Y(_02695_));
 sky130_fd_sc_hd__o31a_1 _05597_ (.A1(_00451_),
    .A2(_00869_),
    .A3(_02156_),
    .B1(_02684_),
    .X(_02706_));
 sky130_fd_sc_hd__nor2_1 _05598_ (.A(_02695_),
    .B(_02706_),
    .Y(_02717_));
 sky130_fd_sc_hd__a22oi_1 _05599_ (.A1(net11),
    .A2(net46),
    .B1(net47),
    .B2(net10),
    .Y(_02728_));
 sky130_fd_sc_hd__and4_1 _05600_ (.A(net11),
    .B(net10),
    .C(net46),
    .D(net47),
    .X(_02739_));
 sky130_fd_sc_hd__o22a_1 _05601_ (.A1(_02728_),
    .A2(_02739_),
    .B1(_00198_),
    .B2(_00781_),
    .X(_02750_));
 sky130_fd_sc_hd__nor4_1 _05602_ (.A(_02728_),
    .B(_00198_),
    .C(_00781_),
    .D(_02739_),
    .Y(_02761_));
 sky130_fd_sc_hd__nor2_1 _05603_ (.A(_02750_),
    .B(_02761_),
    .Y(_02772_));
 sky130_fd_sc_hd__and4_1 _05604_ (.A(net14),
    .B(net13),
    .C(net43),
    .D(net42),
    .X(_02783_));
 sky130_fd_sc_hd__o22a_1 _05605_ (.A1(_00253_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00242_),
    .X(_02794_));
 sky130_fd_sc_hd__and4bb_1 _05606_ (.A_N(_02783_),
    .B_N(_02794_),
    .C(net11),
    .D(net45),
    .X(_02805_));
 sky130_fd_sc_hd__a41o_1 _05607_ (.A1(net14),
    .A2(net13),
    .A3(net43),
    .A4(net42),
    .B1(_02805_),
    .X(_02816_));
 sky130_fd_sc_hd__o2bb2a_1 _05608_ (.A1_N(net13),
    .A2_N(net45),
    .B1(_02178_),
    .B2(_02189_),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_1 _05609_ (.A(_02200_),
    .B(_02827_),
    .Y(_02838_));
 sky130_fd_sc_hd__xor2_1 _05610_ (.A(_02816_),
    .B(_02838_),
    .X(_02849_));
 sky130_fd_sc_hd__or3b_1 _05611_ (.A(_02750_),
    .B(_02761_),
    .C_N(_02849_),
    .X(_02860_));
 sky130_fd_sc_hd__xor2_1 _05612_ (.A(_02772_),
    .B(_02849_),
    .X(_02871_));
 sky130_fd_sc_hd__a21o_1 _05613_ (.A1(_02717_),
    .A2(_02871_),
    .B1(_02695_),
    .X(_02882_));
 sky130_fd_sc_hd__nand2b_1 _05614_ (.A_N(_02167_),
    .B(_02343_),
    .Y(_02893_));
 sky130_fd_sc_hd__nand2_1 _05615_ (.A(_02354_),
    .B(_02893_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2b_1 _05616_ (.A_N(_02904_),
    .B(_02882_),
    .Y(_02915_));
 sky130_fd_sc_hd__o211ai_1 _05617_ (.A1(_02255_),
    .A2(_02310_),
    .B1(_02915_),
    .C1(_02233_),
    .Y(_02926_));
 sky130_fd_sc_hd__a21o_1 _05618_ (.A1(_02233_),
    .A2(_02321_),
    .B1(_02915_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_1 _05619_ (.A(_02926_),
    .B(_02937_),
    .Y(_02948_));
 sky130_fd_sc_hd__xnor2_1 _05620_ (.A(_02618_),
    .B(_02948_),
    .Y(_02959_));
 sky130_fd_sc_hd__or2_1 _05621_ (.A(_02607_),
    .B(_02959_),
    .X(_02970_));
 sky130_fd_sc_hd__o21ai_1 _05622_ (.A1(_02618_),
    .A2(_02948_),
    .B1(_02937_),
    .Y(_02981_));
 sky130_fd_sc_hd__o21ba_1 _05623_ (.A1(_02596_),
    .A2(_02970_),
    .B1_N(_02981_),
    .X(_02992_));
 sky130_fd_sc_hd__xnor2_1 _05624_ (.A(_02596_),
    .B(_02970_),
    .Y(_03003_));
 sky130_fd_sc_hd__a21o_1 _05625_ (.A1(_02596_),
    .A2(_02970_),
    .B1(_02992_),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_1 _05626_ (.A(_02574_),
    .B(_03014_),
    .Y(_03025_));
 sky130_fd_sc_hd__and2_1 _05627_ (.A(_02574_),
    .B(_03014_),
    .X(_03036_));
 sky130_fd_sc_hd__nor2_1 _05628_ (.A(_03025_),
    .B(_03036_),
    .Y(_03047_));
 sky130_fd_sc_hd__a41o_1 _05629_ (.A1(net11),
    .A2(net10),
    .A3(net46),
    .A4(net47),
    .B1(_02761_),
    .X(_03058_));
 sky130_fd_sc_hd__a21bo_1 _05630_ (.A1(_02816_),
    .A2(_02838_),
    .B1_N(_02860_),
    .X(_03069_));
 sky130_fd_sc_hd__o22a_1 _05631_ (.A1(_00242_),
    .A2(_00451_),
    .B1(_02651_),
    .B2(_02662_),
    .X(_03080_));
 sky130_fd_sc_hd__nor2_1 _05632_ (.A(_02673_),
    .B(_03080_),
    .Y(_03091_));
 sky130_fd_sc_hd__and3_1 _05633_ (.A(net14),
    .B(net39),
    .C(_02156_),
    .X(_03102_));
 sky130_fd_sc_hd__a22oi_1 _05634_ (.A1(net15),
    .A2(net39),
    .B1(net40),
    .B2(net14),
    .Y(_03113_));
 sky130_fd_sc_hd__a22o_1 _05635_ (.A1(net15),
    .A2(net39),
    .B1(net40),
    .B2(net14),
    .X(_03124_));
 sky130_fd_sc_hd__and4b_1 _05636_ (.A_N(_03102_),
    .B(_03124_),
    .C(net13),
    .D(net41),
    .X(_03135_));
 sky130_fd_sc_hd__a31o_1 _05637_ (.A1(net13),
    .A2(net41),
    .A3(_03124_),
    .B1(_03102_),
    .X(_03146_));
 sky130_fd_sc_hd__o21ai_1 _05638_ (.A1(_03102_),
    .A2(_03135_),
    .B1(_03091_),
    .Y(_03157_));
 sky130_fd_sc_hd__a311o_1 _05639_ (.A1(net39),
    .A2(_00880_),
    .A3(_02156_),
    .B1(_02640_),
    .C1(_02673_),
    .X(_03168_));
 sky130_fd_sc_hd__and4_1 _05640_ (.A(_02684_),
    .B(_03168_),
    .C(_03091_),
    .D(_03146_),
    .X(_03179_));
 sky130_fd_sc_hd__a22oi_1 _05641_ (.A1(net10),
    .A2(net46),
    .B1(net47),
    .B2(net9),
    .Y(_03190_));
 sky130_fd_sc_hd__and4_1 _05642_ (.A(net9),
    .B(net10),
    .C(net46),
    .D(net47),
    .X(_03201_));
 sky130_fd_sc_hd__a2bb2o_1 _05643_ (.A1_N(_03190_),
    .A2_N(_03201_),
    .B1(net8),
    .B2(net117),
    .X(_03212_));
 sky130_fd_sc_hd__or4_1 _05644_ (.A(_03190_),
    .B(_00209_),
    .C(_00781_),
    .D(_03201_),
    .X(_03223_));
 sky130_fd_sc_hd__and4_1 _05645_ (.A(net11),
    .B(net13),
    .C(net43),
    .D(net42),
    .X(_03234_));
 sky130_fd_sc_hd__or4_1 _05646_ (.A(_00220_),
    .B(_00253_),
    .C(_00462_),
    .D(_00473_),
    .X(_03245_));
 sky130_fd_sc_hd__o22a_1 _05647_ (.A1(_00220_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00253_),
    .X(_03256_));
 sky130_fd_sc_hd__and4b_1 _05648_ (.A_N(_03256_),
    .B(net10),
    .C(_03245_),
    .D(net45),
    .X(_03267_));
 sky130_fd_sc_hd__or4b_1 _05649_ (.A(_00231_),
    .B(_03234_),
    .C(_03256_),
    .D_N(net45),
    .X(_03278_));
 sky130_fd_sc_hd__o2bb2a_1 _05650_ (.A1_N(net11),
    .A2_N(net45),
    .B1(_02783_),
    .B2(_02794_),
    .X(_03289_));
 sky130_fd_sc_hd__o211ai_1 _05651_ (.A1(_02805_),
    .A2(_03289_),
    .B1(_03278_),
    .C1(_03245_),
    .Y(_03300_));
 sky130_fd_sc_hd__a211o_1 _05652_ (.A1(_03245_),
    .A2(_03278_),
    .B1(_03289_),
    .C1(_02805_),
    .X(_03311_));
 sky130_fd_sc_hd__a22o_1 _05653_ (.A1(_03212_),
    .A2(_03223_),
    .B1(_03300_),
    .B2(_03311_),
    .X(_03322_));
 sky130_fd_sc_hd__nand4_1 _05654_ (.A(_03212_),
    .B(_03223_),
    .C(_03300_),
    .D(_03311_),
    .Y(_03333_));
 sky130_fd_sc_hd__a22oi_2 _05655_ (.A1(_03091_),
    .A2(_03146_),
    .B1(_03168_),
    .B2(_02684_),
    .Y(_03344_));
 sky130_fd_sc_hd__nor2_1 _05656_ (.A(_03179_),
    .B(_03344_),
    .Y(_03355_));
 sky130_fd_sc_hd__and3_1 _05657_ (.A(_03355_),
    .B(_03333_),
    .C(_03322_),
    .X(_03366_));
 sky130_fd_sc_hd__xor2_1 _05658_ (.A(_02717_),
    .B(_02871_),
    .X(_03377_));
 sky130_fd_sc_hd__o21a_1 _05659_ (.A1(_03179_),
    .A2(_03366_),
    .B1(_03377_),
    .X(_03388_));
 sky130_fd_sc_hd__o211a_1 _05660_ (.A1(_03179_),
    .A2(_03366_),
    .B1(_03069_),
    .C1(_03377_),
    .X(_03399_));
 sky130_fd_sc_hd__or2_1 _05661_ (.A(_03069_),
    .B(_03388_),
    .X(_03410_));
 sky130_fd_sc_hd__and2b_1 _05662_ (.A_N(_03399_),
    .B(_03410_),
    .X(_03421_));
 sky130_fd_sc_hd__xnor2_1 _05663_ (.A(_03058_),
    .B(_03421_),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2b_1 _05664_ (.A_N(_02882_),
    .B(_02904_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_1 _05665_ (.A(_02915_),
    .B(_03443_),
    .Y(_03454_));
 sky130_fd_sc_hd__or2_1 _05666_ (.A(_03432_),
    .B(_03454_),
    .X(_03465_));
 sky130_fd_sc_hd__nand2_1 _05667_ (.A(_02607_),
    .B(_02959_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _05668_ (.A(_02970_),
    .B(_03476_),
    .Y(_03487_));
 sky130_fd_sc_hd__or3_1 _05669_ (.A(_03432_),
    .B(_03454_),
    .C(_03487_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _05670_ (.A1(_03421_),
    .A2(_03058_),
    .B1(_03399_),
    .X(_03509_));
 sky130_fd_sc_hd__o21ai_1 _05671_ (.A1(_03432_),
    .A2(_03454_),
    .B1(_03487_),
    .Y(_03520_));
 sky130_fd_sc_hd__and2_1 _05672_ (.A(_03498_),
    .B(_03520_),
    .X(_03531_));
 sky130_fd_sc_hd__nand2_1 _05673_ (.A(_03531_),
    .B(_03509_),
    .Y(_03542_));
 sky130_fd_sc_hd__xor2_1 _05674_ (.A(_02981_),
    .B(_03003_),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _05675_ (.A1(_03498_),
    .A2(_03542_),
    .B1(_03553_),
    .Y(_03564_));
 sky130_fd_sc_hd__o211a_1 _05676_ (.A1(_03465_),
    .A2(_03487_),
    .B1(_03542_),
    .C1(_03553_),
    .X(_03575_));
 sky130_fd_sc_hd__nor2_1 _05677_ (.A(_03564_),
    .B(_03575_),
    .Y(_03586_));
 sky130_fd_sc_hd__a211o_1 _05678_ (.A1(_03421_),
    .A2(_03058_),
    .B1(_03399_),
    .C1(_03531_),
    .X(_03597_));
 sky130_fd_sc_hd__nand2_1 _05679_ (.A(_03432_),
    .B(_03454_),
    .Y(_03608_));
 sky130_fd_sc_hd__nand2_1 _05680_ (.A(_03465_),
    .B(_03608_),
    .Y(_03619_));
 sky130_fd_sc_hd__a311oi_1 _05681_ (.A1(_03322_),
    .A2(_03355_),
    .A3(_03333_),
    .B1(_03179_),
    .C1(_03377_),
    .Y(_03630_));
 sky130_fd_sc_hd__or2_1 _05682_ (.A(_03388_),
    .B(_03630_),
    .X(_03641_));
 sky130_fd_sc_hd__nand2b_1 _05683_ (.A_N(_03201_),
    .B(_03223_),
    .Y(_03652_));
 sky130_fd_sc_hd__and2_1 _05684_ (.A(_03311_),
    .B(_03333_),
    .X(_03663_));
 sky130_fd_sc_hd__o2bb2a_1 _05685_ (.A1_N(_03322_),
    .A2_N(_03333_),
    .B1(_03344_),
    .B2(_03179_),
    .X(_03674_));
 sky130_fd_sc_hd__nor2_1 _05686_ (.A(_03366_),
    .B(_03674_),
    .Y(_03685_));
 sky130_fd_sc_hd__and2_2 _05687_ (.A(net15),
    .B(net37),
    .X(_03696_));
 sky130_fd_sc_hd__nand2_1 _05688_ (.A(_00880_),
    .B(net38),
    .Y(_03707_));
 sky130_fd_sc_hd__o22a_1 _05689_ (.A1(_00253_),
    .A2(_00451_),
    .B1(_03102_),
    .B2(_03113_),
    .X(_03718_));
 sky130_fd_sc_hd__nor2_1 _05690_ (.A(_03135_),
    .B(_03718_),
    .Y(_03729_));
 sky130_fd_sc_hd__and4_1 _05691_ (.A(net38),
    .B(_03729_),
    .C(_00880_),
    .D(_03696_),
    .X(_03740_));
 sky130_fd_sc_hd__nand4_2 _05692_ (.A(net14),
    .B(net13),
    .C(net39),
    .D(net40),
    .Y(_03751_));
 sky130_fd_sc_hd__a22o_1 _05693_ (.A1(net14),
    .A2(net39),
    .B1(net40),
    .B2(net13),
    .X(_03762_));
 sky130_fd_sc_hd__nand4_2 _05694_ (.A(_03762_),
    .B(net41),
    .C(net11),
    .D(_03751_),
    .Y(_03773_));
 sky130_fd_sc_hd__a31oi_2 _05695_ (.A1(net38),
    .A2(_00880_),
    .A3(_03696_),
    .B1(_03729_),
    .Y(_03784_));
 sky130_fd_sc_hd__a211oi_2 _05696_ (.A1(_03751_),
    .A2(_03773_),
    .B1(_03784_),
    .C1(_03740_),
    .Y(_03795_));
 sky130_fd_sc_hd__a311o_1 _05697_ (.A1(net13),
    .A2(net41),
    .A3(_03124_),
    .B1(_03102_),
    .C1(_03091_),
    .X(_03806_));
 sky130_fd_sc_hd__o211a_1 _05698_ (.A1(_03740_),
    .A2(_03795_),
    .B1(_03806_),
    .C1(_03157_),
    .X(_03817_));
 sky130_fd_sc_hd__a22oi_2 _05699_ (.A1(net9),
    .A2(net46),
    .B1(net47),
    .B2(net8),
    .Y(_03828_));
 sky130_fd_sc_hd__and4_1 _05700_ (.A(net9),
    .B(net8),
    .C(net46),
    .D(net47),
    .X(_03839_));
 sky130_fd_sc_hd__o22a_1 _05701_ (.A1(_03828_),
    .A2(_03839_),
    .B1(_00176_),
    .B2(_00781_),
    .X(_03850_));
 sky130_fd_sc_hd__nor4_2 _05702_ (.A(_03828_),
    .B(_00176_),
    .C(_00781_),
    .D(_03839_),
    .Y(_03861_));
 sky130_fd_sc_hd__or2_1 _05703_ (.A(_03850_),
    .B(_03861_),
    .X(_03872_));
 sky130_fd_sc_hd__and4_1 _05704_ (.A(net11),
    .B(net10),
    .C(net43),
    .D(net42),
    .X(_03883_));
 sky130_fd_sc_hd__or4_1 _05705_ (.A(_00220_),
    .B(_00231_),
    .C(_00462_),
    .D(_00473_),
    .X(_03894_));
 sky130_fd_sc_hd__o22a_1 _05706_ (.A1(_00231_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00220_),
    .X(_03905_));
 sky130_fd_sc_hd__or4b_2 _05707_ (.A(_00198_),
    .B(_03883_),
    .C(_03905_),
    .D_N(net45),
    .X(_03916_));
 sky130_fd_sc_hd__o2bb2a_1 _05708_ (.A1_N(net10),
    .A2_N(net45),
    .B1(_03234_),
    .B2(_03256_),
    .X(_03927_));
 sky130_fd_sc_hd__o211a_1 _05709_ (.A1(_03267_),
    .A2(_03927_),
    .B1(_03916_),
    .C1(_03894_),
    .X(_03938_));
 sky130_fd_sc_hd__o211ai_1 _05710_ (.A1(_03267_),
    .A2(_03927_),
    .B1(_03916_),
    .C1(_03894_),
    .Y(_03949_));
 sky130_fd_sc_hd__a211o_1 _05711_ (.A1(_03894_),
    .A2(_03916_),
    .B1(_03927_),
    .C1(_03267_),
    .X(_03960_));
 sky130_fd_sc_hd__a2bb2o_1 _05712_ (.A1_N(_03850_),
    .A2_N(_03861_),
    .B1(_03949_),
    .B2(_03960_),
    .X(_03971_));
 sky130_fd_sc_hd__or4b_1 _05713_ (.A(_03850_),
    .B(_03861_),
    .C(_03938_),
    .D_N(_03960_),
    .X(_03982_));
 sky130_fd_sc_hd__and2_1 _05714_ (.A(_03971_),
    .B(_03982_),
    .X(_03993_));
 sky130_fd_sc_hd__a211oi_1 _05715_ (.A1(_03157_),
    .A2(_03806_),
    .B1(_03795_),
    .C1(_03740_),
    .Y(_04004_));
 sky130_fd_sc_hd__nor2_1 _05716_ (.A(_03817_),
    .B(_04004_),
    .Y(_04015_));
 sky130_fd_sc_hd__a21o_1 _05717_ (.A1(_03993_),
    .A2(_04015_),
    .B1(_03817_),
    .X(_04026_));
 sky130_fd_sc_hd__and2_1 _05718_ (.A(_04026_),
    .B(_03685_),
    .X(_04037_));
 sky130_fd_sc_hd__a21boi_1 _05719_ (.A1(_04026_),
    .A2(_03685_),
    .B1_N(_03663_),
    .Y(_04048_));
 sky130_fd_sc_hd__and3b_1 _05720_ (.A_N(_03663_),
    .B(_04026_),
    .C(_03685_),
    .X(_04059_));
 sky130_fd_sc_hd__nor2_1 _05721_ (.A(_04048_),
    .B(_04059_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _05722_ (.A(_03652_),
    .B(_04070_),
    .Y(_04081_));
 sky130_fd_sc_hd__or2_1 _05723_ (.A(_03641_),
    .B(_04081_),
    .X(_04092_));
 sky130_fd_sc_hd__o21ai_1 _05724_ (.A1(_03641_),
    .A2(_04081_),
    .B1(_03619_),
    .Y(_04103_));
 sky130_fd_sc_hd__inv_2 _05725_ (.A(_04103_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _05726_ (.A(_03619_),
    .B(_04092_),
    .Y(_04125_));
 sky130_fd_sc_hd__a21o_1 _05727_ (.A1(_04070_),
    .A2(_03652_),
    .B1(_04059_),
    .X(_04136_));
 sky130_fd_sc_hd__a21o_1 _05728_ (.A1(_04103_),
    .A2(_04136_),
    .B1(_04125_),
    .X(_04147_));
 sky130_fd_sc_hd__and3_1 _05729_ (.A(_03542_),
    .B(_03597_),
    .C(_04147_),
    .X(_04158_));
 sky130_fd_sc_hd__a21oi_1 _05730_ (.A1(_03542_),
    .A2(_03597_),
    .B1(_04147_),
    .Y(_04169_));
 sky130_fd_sc_hd__or2_1 _05731_ (.A(_04158_),
    .B(_04169_),
    .X(_04180_));
 sky130_fd_sc_hd__nand2_1 _05732_ (.A(_03641_),
    .B(_04081_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _05733_ (.A(_04092_),
    .B(_04191_),
    .Y(_04202_));
 sky130_fd_sc_hd__o211a_1 _05734_ (.A1(_03740_),
    .A2(_03784_),
    .B1(_03773_),
    .C1(_03751_),
    .X(_04213_));
 sky130_fd_sc_hd__nor2_1 _05735_ (.A(_03795_),
    .B(_04213_),
    .Y(_04224_));
 sky130_fd_sc_hd__a22o_1 _05736_ (.A1(net11),
    .A2(net41),
    .B1(_03751_),
    .B2(_03762_),
    .X(_04235_));
 sky130_fd_sc_hd__a21oi_1 _05737_ (.A1(_00880_),
    .A2(net36),
    .B1(_03696_),
    .Y(_04246_));
 sky130_fd_sc_hd__and4_1 _05738_ (.A(_00880_),
    .B(net36),
    .C(net37),
    .D(net15),
    .X(_04257_));
 sky130_fd_sc_hd__nand4_1 _05739_ (.A(_00880_),
    .B(net36),
    .C(net37),
    .D(net15),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _05740_ (.A(net14),
    .B(net38),
    .Y(_04279_));
 sky130_fd_sc_hd__o21ai_1 _05741_ (.A1(_04279_),
    .A2(_04246_),
    .B1(_04268_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand3_1 _05742_ (.A(_04290_),
    .B(_04235_),
    .C(_03773_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand4_1 _05743_ (.A(net11),
    .B(net13),
    .C(net39),
    .D(net40),
    .Y(_04312_));
 sky130_fd_sc_hd__a22o_1 _05744_ (.A1(net13),
    .A2(net39),
    .B1(net40),
    .B2(net11),
    .X(_04323_));
 sky130_fd_sc_hd__and4_1 _05745_ (.A(_04323_),
    .B(net41),
    .C(net10),
    .D(_04312_),
    .X(_04334_));
 sky130_fd_sc_hd__a41o_1 _05746_ (.A1(net11),
    .A2(net13),
    .A3(net39),
    .A4(net40),
    .B1(_04334_),
    .X(_04345_));
 sky130_fd_sc_hd__a21o_1 _05747_ (.A1(_03773_),
    .A2(_04235_),
    .B1(_04290_),
    .X(_04356_));
 sky130_fd_sc_hd__and3_1 _05748_ (.A(_04301_),
    .B(_04345_),
    .C(_04356_),
    .X(_04367_));
 sky130_fd_sc_hd__a31o_1 _05749_ (.A1(_03773_),
    .A2(_04235_),
    .A3(_04290_),
    .B1(_04367_),
    .X(_04378_));
 sky130_fd_sc_hd__and2_1 _05750_ (.A(_04224_),
    .B(_04378_),
    .X(_04389_));
 sky130_fd_sc_hd__xnor2_1 _05751_ (.A(_04224_),
    .B(_04378_),
    .Y(_04400_));
 sky130_fd_sc_hd__a22oi_1 _05752_ (.A1(net8),
    .A2(net46),
    .B1(net47),
    .B2(net7),
    .Y(_04411_));
 sky130_fd_sc_hd__and4_1 _05753_ (.A(net7),
    .B(net8),
    .C(net46),
    .D(net47),
    .X(_04422_));
 sky130_fd_sc_hd__a2bb2o_1 _05754_ (.A1_N(_04411_),
    .A2_N(_04422_),
    .B1(net6),
    .B2(net117),
    .X(_04433_));
 sky130_fd_sc_hd__or4_1 _05755_ (.A(_04411_),
    .B(_00187_),
    .C(_00781_),
    .D(_04422_),
    .X(_04444_));
 sky130_fd_sc_hd__nand2_1 _05756_ (.A(_04433_),
    .B(_04444_),
    .Y(_04455_));
 sky130_fd_sc_hd__and4_1 _05757_ (.A(net9),
    .B(net10),
    .C(net43),
    .D(net42),
    .X(_04466_));
 sky130_fd_sc_hd__o22a_1 _05758_ (.A1(_00198_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00231_),
    .X(_04477_));
 sky130_fd_sc_hd__and4bb_1 _05759_ (.A_N(_04466_),
    .B_N(_04477_),
    .C(net8),
    .D(net45),
    .X(_04488_));
 sky130_fd_sc_hd__a41o_1 _05760_ (.A1(net9),
    .A2(net10),
    .A3(net43),
    .A4(net42),
    .B1(_04488_),
    .X(_04499_));
 sky130_fd_sc_hd__a2bb2o_1 _05761_ (.A1_N(_03883_),
    .A2_N(_03905_),
    .B1(net9),
    .B2(net45),
    .X(_04510_));
 sky130_fd_sc_hd__a21oi_1 _05762_ (.A1(_03916_),
    .A2(_04510_),
    .B1(_04499_),
    .Y(_04521_));
 sky130_fd_sc_hd__and3_1 _05763_ (.A(_03916_),
    .B(_04499_),
    .C(_04510_),
    .X(_04532_));
 sky130_fd_sc_hd__nor2_1 _05764_ (.A(_04521_),
    .B(_04532_),
    .Y(_04543_));
 sky130_fd_sc_hd__xor2_1 _05765_ (.A(_04455_),
    .B(_04543_),
    .X(_04554_));
 sky130_fd_sc_hd__nor2_1 _05766_ (.A(_04400_),
    .B(_04554_),
    .Y(_04565_));
 sky130_fd_sc_hd__xor2_1 _05767_ (.A(_03993_),
    .B(_04015_),
    .X(_04576_));
 sky130_fd_sc_hd__o21ai_2 _05768_ (.A1(_04389_),
    .A2(_04565_),
    .B1(_04576_),
    .Y(_04587_));
 sky130_fd_sc_hd__a21o_1 _05769_ (.A1(_03960_),
    .A2(_03982_),
    .B1(_04587_),
    .X(_04598_));
 sky130_fd_sc_hd__o211ai_2 _05770_ (.A1(_03872_),
    .A2(_03938_),
    .B1(_03960_),
    .C1(_04587_),
    .Y(_04609_));
 sky130_fd_sc_hd__o211ai_2 _05771_ (.A1(_03839_),
    .A2(_03861_),
    .B1(_04598_),
    .C1(_04609_),
    .Y(_04620_));
 sky130_fd_sc_hd__inv_2 _05772_ (.A(_04620_),
    .Y(_04631_));
 sky130_fd_sc_hd__a211oi_1 _05773_ (.A1(_04598_),
    .A2(_04609_),
    .B1(_03839_),
    .C1(_03861_),
    .Y(_04641_));
 sky130_fd_sc_hd__nor2_1 _05774_ (.A(_03685_),
    .B(_04026_),
    .Y(_04651_));
 sky130_fd_sc_hd__or2_1 _05775_ (.A(_04037_),
    .B(_04651_),
    .X(_04661_));
 sky130_fd_sc_hd__or3_2 _05776_ (.A(_04661_),
    .B(_04641_),
    .C(_04631_),
    .X(_04671_));
 sky130_fd_sc_hd__or4_1 _05777_ (.A(_04631_),
    .B(_04641_),
    .C(_04661_),
    .D(_04202_),
    .X(_04680_));
 sky130_fd_sc_hd__nand2_1 _05778_ (.A(_04202_),
    .B(_04671_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_1 _05779_ (.A(_04680_),
    .B(_04690_),
    .Y(_04700_));
 sky130_fd_sc_hd__a21o_1 _05780_ (.A1(_04598_),
    .A2(_04620_),
    .B1(_04700_),
    .X(_04709_));
 sky130_fd_sc_hd__inv_2 _05781_ (.A(_04709_),
    .Y(_04719_));
 sky130_fd_sc_hd__o21ai_1 _05782_ (.A1(_04114_),
    .A2(_04125_),
    .B1(_04136_),
    .Y(_04729_));
 sky130_fd_sc_hd__or3_1 _05783_ (.A(_04136_),
    .B(_04125_),
    .C(_04114_),
    .X(_04738_));
 sky130_fd_sc_hd__and2_1 _05784_ (.A(_04729_),
    .B(_04738_),
    .X(_04748_));
 sky130_fd_sc_hd__a21oi_1 _05785_ (.A1(_04680_),
    .A2(_04709_),
    .B1(_04748_),
    .Y(_04758_));
 sky130_fd_sc_hd__o211a_1 _05786_ (.A1(_04202_),
    .A2(_04671_),
    .B1(_04709_),
    .C1(_04748_),
    .X(_04767_));
 sky130_fd_sc_hd__or2_1 _05787_ (.A(_04758_),
    .B(_04767_),
    .X(_04777_));
 sky130_fd_sc_hd__inv_2 _05788_ (.A(_04777_),
    .Y(_04786_));
 sky130_fd_sc_hd__and3_1 _05789_ (.A(_04598_),
    .B(_04620_),
    .C(_04700_),
    .X(_04796_));
 sky130_fd_sc_hd__nor2_1 _05790_ (.A(_04719_),
    .B(_04796_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_1 _05791_ (.A1(_04631_),
    .A2(_04641_),
    .B1(_04661_),
    .Y(_04816_));
 sky130_fd_sc_hd__or3_1 _05792_ (.A(_04389_),
    .B(_04565_),
    .C(_04576_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2_1 _05793_ (.A(_04587_),
    .B(_04826_),
    .Y(_04836_));
 sky130_fd_sc_hd__and4_1 _05794_ (.A(net14),
    .B(net15),
    .C(net37),
    .D(net36),
    .X(_04846_));
 sky130_fd_sc_hd__a22oi_1 _05795_ (.A1(net14),
    .A2(net37),
    .B1(net36),
    .B2(net15),
    .Y(_04856_));
 sky130_fd_sc_hd__and4bb_1 _05796_ (.A_N(_04846_),
    .B_N(_04856_),
    .C(net13),
    .D(net38),
    .X(_04866_));
 sky130_fd_sc_hd__nor2_1 _05797_ (.A(_04846_),
    .B(_04866_),
    .Y(_04877_));
 sky130_fd_sc_hd__o2bb2a_1 _05798_ (.A1_N(_04312_),
    .A2_N(_04323_),
    .B1(_00231_),
    .B2(_00451_),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _05799_ (.A(_04334_),
    .B(_04887_),
    .Y(_04896_));
 sky130_fd_sc_hd__or3_1 _05800_ (.A(_04334_),
    .B(_04877_),
    .C(_04887_),
    .X(_04898_));
 sky130_fd_sc_hd__nand4_2 _05801_ (.A(net11),
    .B(net10),
    .C(net39),
    .D(net40),
    .Y(_04899_));
 sky130_fd_sc_hd__a22o_1 _05802_ (.A1(net11),
    .A2(net39),
    .B1(net40),
    .B2(net10),
    .X(_04900_));
 sky130_fd_sc_hd__nand4_2 _05803_ (.A(_04900_),
    .B(net41),
    .C(net9),
    .D(_04899_),
    .Y(_04901_));
 sky130_fd_sc_hd__nand2_1 _05804_ (.A(_04899_),
    .B(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__xnor2_1 _05805_ (.A(_04877_),
    .B(_04896_),
    .Y(_04903_));
 sky130_fd_sc_hd__a21bo_1 _05806_ (.A1(_04902_),
    .A2(_04903_),
    .B1_N(_04898_),
    .X(_04904_));
 sky130_fd_sc_hd__a21oi_1 _05807_ (.A1(_04301_),
    .A2(_04356_),
    .B1(_04345_),
    .Y(_04905_));
 sky130_fd_sc_hd__nor2_1 _05808_ (.A(_04367_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2_1 _05809_ (.A(_04906_),
    .B(_04904_),
    .Y(_04907_));
 sky130_fd_sc_hd__xnor2_2 _05810_ (.A(_04904_),
    .B(_04906_),
    .Y(_04908_));
 sky130_fd_sc_hd__a22oi_1 _05811_ (.A1(net7),
    .A2(net46),
    .B1(net47),
    .B2(net6),
    .Y(_04909_));
 sky130_fd_sc_hd__and4_1 _05812_ (.A(net7),
    .B(net6),
    .C(net46),
    .D(net47),
    .X(_04910_));
 sky130_fd_sc_hd__o22a_1 _05813_ (.A1(_04909_),
    .A2(_04910_),
    .B1(_00154_),
    .B2(_00781_),
    .X(_04911_));
 sky130_fd_sc_hd__nor4_1 _05814_ (.A(_04909_),
    .B(_00154_),
    .C(_00781_),
    .D(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__and4_1 _05815_ (.A(net9),
    .B(net8),
    .C(net43),
    .D(net42),
    .X(_04913_));
 sky130_fd_sc_hd__o22a_1 _05816_ (.A1(_00209_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00198_),
    .X(_04914_));
 sky130_fd_sc_hd__and4bb_1 _05817_ (.A_N(_04913_),
    .B_N(_04914_),
    .C(net7),
    .D(net45),
    .X(_04915_));
 sky130_fd_sc_hd__a41o_1 _05818_ (.A1(net9),
    .A2(net8),
    .A3(net43),
    .A4(net42),
    .B1(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__o2bb2a_1 _05819_ (.A1_N(net8),
    .A2_N(net45),
    .B1(_04466_),
    .B2(_04477_),
    .X(_04917_));
 sky130_fd_sc_hd__nor2_1 _05820_ (.A(_04488_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__nor2_1 _05821_ (.A(_04918_),
    .B(_04916_),
    .Y(_04919_));
 sky130_fd_sc_hd__o21a_1 _05822_ (.A1(_04913_),
    .A2(_04915_),
    .B1(_04918_),
    .X(_04920_));
 sky130_fd_sc_hd__or2_1 _05823_ (.A(_04919_),
    .B(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__nor3_1 _05824_ (.A(_04911_),
    .B(_04912_),
    .C(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21a_1 _05825_ (.A1(_04911_),
    .A2(_04912_),
    .B1(_04921_),
    .X(_04923_));
 sky130_fd_sc_hd__or2_1 _05826_ (.A(_04922_),
    .B(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__o21ai_1 _05827_ (.A1(_04908_),
    .A2(_04924_),
    .B1(_04907_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand2_1 _05828_ (.A(_04400_),
    .B(_04554_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2b_1 _05829_ (.A_N(_04565_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2b_1 _05830_ (.A_N(_04925_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2b_1 _05831_ (.A_N(_04927_),
    .B(_04925_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _05832_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nor3_1 _05833_ (.A(_03707_),
    .B(_04836_),
    .C(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__o21ai_1 _05834_ (.A1(_03707_),
    .A2(_04930_),
    .B1(_04836_),
    .Y(_04932_));
 sky130_fd_sc_hd__nand2b_1 _05835_ (.A_N(_04931_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2b_1 _05836_ (.A_N(_04422_),
    .B(_04444_),
    .Y(_04934_));
 sky130_fd_sc_hd__a31oi_1 _05837_ (.A1(_04543_),
    .A2(_04444_),
    .A3(_04433_),
    .B1(_04532_),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _05838_ (.A(_04929_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__or3b_1 _05839_ (.A(_04927_),
    .B(_04935_),
    .C_N(_04925_),
    .X(_04937_));
 sky130_fd_sc_hd__a21oi_1 _05840_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04934_),
    .Y(_04938_));
 sky130_fd_sc_hd__and3_1 _05841_ (.A(_04934_),
    .B(_04936_),
    .C(_04937_),
    .X(_04939_));
 sky130_fd_sc_hd__nor2_1 _05842_ (.A(_04938_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__and3b_1 _05843_ (.A_N(_04931_),
    .B(_04940_),
    .C(_04932_),
    .X(_04941_));
 sky130_fd_sc_hd__o211a_1 _05844_ (.A1(_04931_),
    .A2(_04941_),
    .B1(_04671_),
    .C1(_04816_),
    .X(_04942_));
 sky130_fd_sc_hd__a211oi_1 _05845_ (.A1(_04671_),
    .A2(_04816_),
    .B1(_04931_),
    .C1(_04941_),
    .Y(_04943_));
 sky130_fd_sc_hd__or2_1 _05846_ (.A(_04942_),
    .B(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__a21boi_1 _05847_ (.A1(_04934_),
    .A2(_04936_),
    .B1_N(_04937_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ba_2 _05848_ (.A1(_04943_),
    .A2(_04945_),
    .B1_N(_04942_),
    .X(_04946_));
 sky130_fd_sc_hd__xor2_1 _05849_ (.A(_04944_),
    .B(_04945_),
    .X(_04947_));
 sky130_fd_sc_hd__xnor2_2 _05850_ (.A(_04933_),
    .B(_04940_),
    .Y(_04948_));
 sky130_fd_sc_hd__xor2_1 _05851_ (.A(_03707_),
    .B(_04930_),
    .X(_04949_));
 sky130_fd_sc_hd__a22oi_2 _05852_ (.A1(net15),
    .A2(net38),
    .B1(_00880_),
    .B2(net37),
    .Y(_04950_));
 sky130_fd_sc_hd__a31oi_4 _05853_ (.A1(net38),
    .A2(_00880_),
    .A3(_03696_),
    .B1(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__and4_1 _05854_ (.A(net14),
    .B(net13),
    .C(net37),
    .D(net36),
    .X(_04952_));
 sky130_fd_sc_hd__nand2_1 _05855_ (.A(net11),
    .B(net38),
    .Y(_04953_));
 sky130_fd_sc_hd__a22oi_2 _05856_ (.A1(net13),
    .A2(net37),
    .B1(net36),
    .B2(net14),
    .Y(_04954_));
 sky130_fd_sc_hd__nor3_1 _05857_ (.A(_04953_),
    .B(_04954_),
    .C(_04952_),
    .Y(_04955_));
 sky130_fd_sc_hd__o21bai_1 _05858_ (.A1(_04953_),
    .A2(_04954_),
    .B1_N(_04952_),
    .Y(_04956_));
 sky130_fd_sc_hd__a22o_1 _05859_ (.A1(net9),
    .A2(net41),
    .B1(_04899_),
    .B2(_04900_),
    .X(_04957_));
 sky130_fd_sc_hd__o211ai_2 _05860_ (.A1(_04952_),
    .A2(_04955_),
    .B1(_04957_),
    .C1(_04901_),
    .Y(_04958_));
 sky130_fd_sc_hd__nand4_1 _05861_ (.A(net9),
    .B(net10),
    .C(net39),
    .D(net40),
    .Y(_04959_));
 sky130_fd_sc_hd__a22o_1 _05862_ (.A1(net10),
    .A2(net39),
    .B1(net40),
    .B2(net9),
    .X(_04960_));
 sky130_fd_sc_hd__nand4_1 _05863_ (.A(_04960_),
    .B(net41),
    .C(net8),
    .D(_04959_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand2_1 _05864_ (.A(_04959_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__a21o_1 _05865_ (.A1(_04901_),
    .A2(_04957_),
    .B1(_04956_),
    .X(_04963_));
 sky130_fd_sc_hd__and3_1 _05866_ (.A(_04958_),
    .B(_04962_),
    .C(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__nand3_1 _05867_ (.A(_04958_),
    .B(_04962_),
    .C(_04963_),
    .Y(_04965_));
 sky130_fd_sc_hd__a31o_1 _05868_ (.A1(_04901_),
    .A2(_04956_),
    .A3(_04957_),
    .B1(_04964_),
    .X(_04966_));
 sky130_fd_sc_hd__xor2_1 _05869_ (.A(_04902_),
    .B(_04903_),
    .X(_04967_));
 sky130_fd_sc_hd__a22oi_2 _05870_ (.A1(net6),
    .A2(net46),
    .B1(net47),
    .B2(net5),
    .Y(_04968_));
 sky130_fd_sc_hd__and4_1 _05871_ (.A(net5),
    .B(net6),
    .C(net46),
    .D(net47),
    .X(_04969_));
 sky130_fd_sc_hd__o22a_1 _05872_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_00165_),
    .B2(_00781_),
    .X(_04970_));
 sky130_fd_sc_hd__nor4_2 _05873_ (.A(_04968_),
    .B(_00165_),
    .C(_00781_),
    .D(_04969_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand4_4 _05874_ (.A(net7),
    .B(net8),
    .C(net43),
    .D(net42),
    .Y(_04972_));
 sky130_fd_sc_hd__a22o_1 _05875_ (.A1(net7),
    .A2(net43),
    .B1(net42),
    .B2(net8),
    .X(_04973_));
 sky130_fd_sc_hd__nand4_4 _05876_ (.A(_04973_),
    .B(net45),
    .C(net6),
    .D(_04972_),
    .Y(_04974_));
 sky130_fd_sc_hd__o2bb2a_1 _05877_ (.A1_N(net7),
    .A2_N(net45),
    .B1(_04913_),
    .B2(_04914_),
    .X(_04975_));
 sky130_fd_sc_hd__a211o_1 _05878_ (.A1(_04972_),
    .A2(_04974_),
    .B1(_04975_),
    .C1(_04915_),
    .X(_04976_));
 sky130_fd_sc_hd__o211ai_1 _05879_ (.A1(_04915_),
    .A2(_04975_),
    .B1(_04974_),
    .C1(_04972_),
    .Y(_04977_));
 sky130_fd_sc_hd__or4bb_2 _05880_ (.A(_04970_),
    .B(_04971_),
    .C_N(_04976_),
    .D_N(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__a2bb2o_1 _05881_ (.A1_N(_04970_),
    .A2_N(_04971_),
    .B1(_04976_),
    .B2(_04977_),
    .X(_04979_));
 sky130_fd_sc_hd__nand2_1 _05882_ (.A(_04978_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__xnor2_1 _05883_ (.A(_04966_),
    .B(_04967_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _05884_ (.A(_04980_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__a21o_1 _05885_ (.A1(_04966_),
    .A2(_04967_),
    .B1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__nor2_2 _05886_ (.A(_00264_),
    .B(_00418_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_2 _05887_ (.A(net15),
    .B(net34),
    .Y(_04985_));
 sky130_fd_sc_hd__o2bb2a_1 _05888_ (.A1_N(net13),
    .A2_N(net38),
    .B1(_04846_),
    .B2(_04856_),
    .X(_04986_));
 sky130_fd_sc_hd__nor2_1 _05889_ (.A(_04866_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__and4_1 _05890_ (.A(net116),
    .B(_04987_),
    .C(_04985_),
    .D(net35),
    .X(_04988_));
 sky130_fd_sc_hd__o2bb2a_1 _05891_ (.A1_N(net14),
    .A2_N(net38),
    .B1(_04246_),
    .B2(_04257_),
    .X(_04989_));
 sky130_fd_sc_hd__and4b_1 _05892_ (.A_N(_04246_),
    .B(_04268_),
    .C(net14),
    .D(net38),
    .X(_04990_));
 sky130_fd_sc_hd__nor2_1 _05893_ (.A(_04989_),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__o2111ai_4 _05894_ (.A1(_04984_),
    .A2(_04987_),
    .B1(_00880_),
    .C1(_04991_),
    .D1(net35),
    .Y(_04992_));
 sky130_fd_sc_hd__xnor2_2 _05895_ (.A(_04908_),
    .B(_04924_),
    .Y(_04993_));
 sky130_fd_sc_hd__nor2_1 _05896_ (.A(_04992_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__xor2_2 _05897_ (.A(_04992_),
    .B(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__xor2_2 _05898_ (.A(_04983_),
    .B(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__nand3_1 _05899_ (.A(_04949_),
    .B(_04951_),
    .C(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a21o_1 _05900_ (.A1(_04951_),
    .A2(_04996_),
    .B1(_04949_),
    .X(_04998_));
 sky130_fd_sc_hd__and2_1 _05901_ (.A(_04997_),
    .B(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__a41o_1 _05902_ (.A1(net7),
    .A2(net6),
    .A3(net46),
    .A4(net47),
    .B1(_04912_),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_1 _05903_ (.A1(_04995_),
    .A2(_04983_),
    .B1(_04994_),
    .X(_05001_));
 sky130_fd_sc_hd__o21a_1 _05904_ (.A1(_04920_),
    .A2(_04922_),
    .B1(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__a211oi_1 _05905_ (.A1(_04916_),
    .A2(_04918_),
    .B1(_04922_),
    .C1(_05001_),
    .Y(_05003_));
 sky130_fd_sc_hd__nor2_1 _05906_ (.A(_05002_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__xor2_1 _05907_ (.A(_05000_),
    .B(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__a21bo_1 _05908_ (.A1(_05005_),
    .A2(_04998_),
    .B1_N(_04997_),
    .X(_05006_));
 sky130_fd_sc_hd__nand2_1 _05909_ (.A(_05006_),
    .B(_04948_),
    .Y(_05007_));
 sky130_fd_sc_hd__xnor2_2 _05910_ (.A(_04948_),
    .B(_05006_),
    .Y(_05008_));
 sky130_fd_sc_hd__a21oi_2 _05911_ (.A1(_05004_),
    .A2(_05000_),
    .B1(_05002_),
    .Y(_05009_));
 sky130_fd_sc_hd__o21ai_1 _05912_ (.A1(_05009_),
    .A2(_05008_),
    .B1(_05007_),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_1 _05913_ (.A(_05010_),
    .B(_04947_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _05914_ (.A(_04947_),
    .B(_05010_),
    .Y(_05012_));
 sky130_fd_sc_hd__and2b_1 _05915_ (.A_N(_05011_),
    .B(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__xnor2_2 _05916_ (.A(_05008_),
    .B(_05009_),
    .Y(_05014_));
 sky130_fd_sc_hd__a311o_1 _05917_ (.A1(net35),
    .A2(_00880_),
    .A3(_04984_),
    .B1(_04988_),
    .C1(_04991_),
    .X(_05015_));
 sky130_fd_sc_hd__nand2_1 _05918_ (.A(_04992_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__and4_1 _05919_ (.A(net11),
    .B(net13),
    .C(net37),
    .D(net36),
    .X(_05017_));
 sky130_fd_sc_hd__o2bb2a_1 _05920_ (.A1_N(net11),
    .A2_N(net37),
    .B1(_00429_),
    .B2(_00253_),
    .X(_05018_));
 sky130_fd_sc_hd__a22o_1 _05921_ (.A1(net11),
    .A2(net37),
    .B1(net36),
    .B2(net13),
    .X(_05019_));
 sky130_fd_sc_hd__and4b_1 _05922_ (.A_N(_05017_),
    .B(_05019_),
    .C(net10),
    .D(net38),
    .X(_05020_));
 sky130_fd_sc_hd__a31o_1 _05923_ (.A1(_05019_),
    .A2(net38),
    .A3(net10),
    .B1(_05017_),
    .X(_05021_));
 sky130_fd_sc_hd__a22o_1 _05924_ (.A1(net8),
    .A2(net41),
    .B1(_04959_),
    .B2(_04960_),
    .X(_05022_));
 sky130_fd_sc_hd__nand3_1 _05925_ (.A(_04961_),
    .B(_05021_),
    .C(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand4_2 _05926_ (.A(net9),
    .B(net8),
    .C(net39),
    .D(net40),
    .Y(_05024_));
 sky130_fd_sc_hd__a22o_1 _05927_ (.A1(net9),
    .A2(net39),
    .B1(net40),
    .B2(net8),
    .X(_05025_));
 sky130_fd_sc_hd__nand4_2 _05928_ (.A(_05025_),
    .B(net41),
    .C(net7),
    .D(_05024_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _05929_ (.A(_05024_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__a21o_1 _05930_ (.A1(_04961_),
    .A2(_05022_),
    .B1(_05021_),
    .X(_05028_));
 sky130_fd_sc_hd__a21boi_2 _05931_ (.A1(_05027_),
    .A2(_05028_),
    .B1_N(_05023_),
    .Y(_05029_));
 sky130_fd_sc_hd__a21o_1 _05932_ (.A1(_04958_),
    .A2(_04963_),
    .B1(_04962_),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_1 _05933_ (.A(_04965_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__or3b_1 _05934_ (.A(_04964_),
    .B(_05029_),
    .C_N(_05030_),
    .X(_05032_));
 sky130_fd_sc_hd__xnor2_1 _05935_ (.A(_05029_),
    .B(_05031_),
    .Y(_05033_));
 sky130_fd_sc_hd__and4_1 _05936_ (.A(net5),
    .B(net4),
    .C(net46),
    .D(net47),
    .X(_05034_));
 sky130_fd_sc_hd__a22oi_1 _05937_ (.A1(net5),
    .A2(net46),
    .B1(net47),
    .B2(net4),
    .Y(_05035_));
 sky130_fd_sc_hd__a22o_1 _05938_ (.A1(net5),
    .A2(net46),
    .B1(net47),
    .B2(net4),
    .X(_05036_));
 sky130_fd_sc_hd__and4b_1 _05939_ (.A_N(_05034_),
    .B(net3),
    .C(net117),
    .D(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__o22a_1 _05940_ (.A1(_05034_),
    .A2(_05035_),
    .B1(_00132_),
    .B2(_00781_),
    .X(_05038_));
 sky130_fd_sc_hd__or2_1 _05941_ (.A(_05037_),
    .B(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__nand4_1 _05942_ (.A(net7),
    .B(net6),
    .C(net43),
    .D(net42),
    .Y(_05040_));
 sky130_fd_sc_hd__a22o_1 _05943_ (.A1(net6),
    .A2(net43),
    .B1(net42),
    .B2(net7),
    .X(_05041_));
 sky130_fd_sc_hd__nand4_1 _05944_ (.A(_05041_),
    .B(net45),
    .C(net5),
    .D(_05040_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _05945_ (.A(_05040_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__a22o_1 _05946_ (.A1(net6),
    .A2(net45),
    .B1(_04972_),
    .B2(_04973_),
    .X(_05044_));
 sky130_fd_sc_hd__nand3_1 _05947_ (.A(_04974_),
    .B(_05043_),
    .C(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a21o_1 _05948_ (.A1(_04974_),
    .A2(_05044_),
    .B1(_05043_),
    .X(_05046_));
 sky130_fd_sc_hd__nand2_1 _05949_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nor2_1 _05950_ (.A(_05039_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__o21ai_1 _05951_ (.A1(_05037_),
    .A2(_05038_),
    .B1(_05047_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2b_1 _05952_ (.A_N(_05048_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__or2_1 _05953_ (.A(_05033_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o32a_1 _05954_ (.A1(_04984_),
    .A2(_00407_),
    .A3(_00869_),
    .B1(_04986_),
    .B2(_04866_),
    .X(_05052_));
 sky130_fd_sc_hd__nor2_1 _05955_ (.A(_04988_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__o22a_1 _05956_ (.A1(_00264_),
    .A2(_00407_),
    .B1(_00418_),
    .B2(_00869_),
    .X(_05054_));
 sky130_fd_sc_hd__a31oi_1 _05957_ (.A1(net35),
    .A2(net116),
    .A3(_04984_),
    .B1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _05958_ (.A(net15),
    .B(net64),
    .Y(_05056_));
 sky130_fd_sc_hd__nand4_2 _05959_ (.A(net116),
    .B(net34),
    .C(net64),
    .D(net15),
    .Y(_05057_));
 sky130_fd_sc_hd__a22o_1 _05960_ (.A1(net15),
    .A2(net34),
    .B1(net116),
    .B2(net64),
    .X(_05058_));
 sky130_fd_sc_hd__and4_1 _05961_ (.A(_05058_),
    .B(net35),
    .C(net14),
    .D(_05057_),
    .X(_05059_));
 sky130_fd_sc_hd__nand4_2 _05962_ (.A(_05058_),
    .B(net35),
    .C(net14),
    .D(_05057_),
    .Y(_05060_));
 sky130_fd_sc_hd__a311o_1 _05963_ (.A1(net64),
    .A2(net116),
    .A3(_04984_),
    .B1(_05055_),
    .C1(_05059_),
    .X(_05061_));
 sky130_fd_sc_hd__a21bo_1 _05964_ (.A1(_05057_),
    .A2(_05060_),
    .B1_N(_05055_),
    .X(_05062_));
 sky130_fd_sc_hd__o2bb2a_1 _05965_ (.A1_N(net11),
    .A2_N(net38),
    .B1(_04952_),
    .B2(_04954_),
    .X(_05063_));
 sky130_fd_sc_hd__nor2_1 _05966_ (.A(_04955_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__a21bo_1 _05967_ (.A1(_05061_),
    .A2(_05064_),
    .B1_N(_05062_),
    .X(_05065_));
 sky130_fd_sc_hd__nand2_2 _05968_ (.A(_05053_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__xnor2_1 _05969_ (.A(_04980_),
    .B(_04981_),
    .Y(_05067_));
 sky130_fd_sc_hd__or2_1 _05970_ (.A(_05066_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _05971_ (.A(_05066_),
    .B(_05067_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_1 _05972_ (.A(_05068_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__a21o_1 _05973_ (.A1(_05032_),
    .A2(_05051_),
    .B1(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__o211ai_1 _05974_ (.A1(_05029_),
    .A2(_05031_),
    .B1(_05051_),
    .C1(_05070_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _05975_ (.A(_05071_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__or2_1 _05976_ (.A(_05016_),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__xnor2_1 _05977_ (.A(_04951_),
    .B(_04996_),
    .Y(_05075_));
 sky130_fd_sc_hd__or3_1 _05978_ (.A(_05016_),
    .B(_05073_),
    .C(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__nand2_1 _05979_ (.A(_04976_),
    .B(_04978_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21ai_1 _05980_ (.A1(_05066_),
    .A2(_05067_),
    .B1(_05071_),
    .Y(_05078_));
 sky130_fd_sc_hd__a22oi_2 _05981_ (.A1(_04976_),
    .A2(_04978_),
    .B1(_05068_),
    .B2(_05071_),
    .Y(_05079_));
 sky130_fd_sc_hd__o2111ai_1 _05982_ (.A1(_05066_),
    .A2(_05067_),
    .B1(_05071_),
    .C1(_04978_),
    .D1(_04976_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand2b_1 _05983_ (.A_N(_05079_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__o21ba_1 _05984_ (.A1(_04969_),
    .A2(_04971_),
    .B1_N(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__o21a_1 _05985_ (.A1(_04969_),
    .A2(_04971_),
    .B1(_05081_),
    .X(_05083_));
 sky130_fd_sc_hd__nor3_1 _05986_ (.A(_04969_),
    .B(_04971_),
    .C(_05081_),
    .Y(_05084_));
 sky130_fd_sc_hd__nor2_1 _05987_ (.A(_05083_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__xnor2_1 _05988_ (.A(_05074_),
    .B(_05075_),
    .Y(_05086_));
 sky130_fd_sc_hd__or2_1 _05989_ (.A(_05085_),
    .B(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__xnor2_1 _05990_ (.A(_04999_),
    .B(_05005_),
    .Y(_05088_));
 sky130_fd_sc_hd__a21o_1 _05991_ (.A1(_05076_),
    .A2(_05087_),
    .B1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__o211ai_1 _05992_ (.A1(_05074_),
    .A2(_05075_),
    .B1(_05087_),
    .C1(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__and2_1 _05993_ (.A(_05089_),
    .B(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__o21a_1 _05994_ (.A1(_05079_),
    .A2(_05082_),
    .B1(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__o21ai_1 _05995_ (.A1(_05079_),
    .A2(_05082_),
    .B1(_05091_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _05996_ (.A(_05089_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__a21o_1 _05997_ (.A1(_05089_),
    .A2(_05093_),
    .B1(_05014_),
    .X(_05095_));
 sky130_fd_sc_hd__xnor2_2 _05998_ (.A(_05014_),
    .B(_05094_),
    .Y(_05096_));
 sky130_fd_sc_hd__a211oi_1 _05999_ (.A1(_05077_),
    .A2(_05078_),
    .B1(_05082_),
    .C1(_05091_),
    .Y(_05097_));
 sky130_fd_sc_hd__nor2_1 _06000_ (.A(_05092_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__and4_1 _06001_ (.A(net11),
    .B(net10),
    .C(net37),
    .D(net36),
    .X(_05099_));
 sky130_fd_sc_hd__a22oi_1 _06002_ (.A1(net10),
    .A2(net37),
    .B1(net36),
    .B2(net11),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _06003_ (.A(net9),
    .B(net38),
    .Y(_05101_));
 sky130_fd_sc_hd__or3_1 _06004_ (.A(_05101_),
    .B(_05100_),
    .C(_05099_),
    .X(_05102_));
 sky130_fd_sc_hd__o21bai_1 _06005_ (.A1(_05100_),
    .A2(_05101_),
    .B1_N(_05099_),
    .Y(_05103_));
 sky130_fd_sc_hd__a22o_1 _06006_ (.A1(net7),
    .A2(net41),
    .B1(_05024_),
    .B2(_05025_),
    .X(_05104_));
 sky130_fd_sc_hd__nand3_1 _06007_ (.A(_05026_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2_1 _06008_ (.A(net7),
    .B(net39),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_1 _06009_ (.A(net7),
    .B(net40),
    .Y(_05107_));
 sky130_fd_sc_hd__and4_1 _06010_ (.A(net7),
    .B(net8),
    .C(net39),
    .D(net40),
    .X(_05108_));
 sky130_fd_sc_hd__a22oi_1 _06011_ (.A1(net8),
    .A2(net39),
    .B1(net40),
    .B2(net7),
    .Y(_05109_));
 sky130_fd_sc_hd__a22o_1 _06012_ (.A1(net8),
    .A2(net39),
    .B1(net40),
    .B2(net7),
    .X(_05110_));
 sky130_fd_sc_hd__nor4_1 _06013_ (.A(_00187_),
    .B(_05109_),
    .C(_00451_),
    .D(_05108_),
    .Y(_05111_));
 sky130_fd_sc_hd__a31o_1 _06014_ (.A1(_05110_),
    .A2(net41),
    .A3(net6),
    .B1(_05108_),
    .X(_05112_));
 sky130_fd_sc_hd__a21o_1 _06015_ (.A1(_05026_),
    .A2(_05104_),
    .B1(_05103_),
    .X(_05113_));
 sky130_fd_sc_hd__and3_1 _06016_ (.A(_05105_),
    .B(_05112_),
    .C(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__a21boi_1 _06017_ (.A1(_05112_),
    .A2(_05113_),
    .B1_N(_05105_),
    .Y(_05115_));
 sky130_fd_sc_hd__a22o_1 _06018_ (.A1(_05024_),
    .A2(_05026_),
    .B1(_05028_),
    .B2(_05023_),
    .X(_05116_));
 sky130_fd_sc_hd__nand3b_1 _06019_ (.A_N(_05027_),
    .B(_05028_),
    .C(_05023_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _06020_ (.A(_05116_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__a21o_1 _06021_ (.A1(_05116_),
    .A2(_05117_),
    .B1(_05115_),
    .X(_05119_));
 sky130_fd_sc_hd__xor2_1 _06022_ (.A(_05115_),
    .B(_05118_),
    .X(_05120_));
 sky130_fd_sc_hd__or4b_2 _06023_ (.A(_00132_),
    .B(_00165_),
    .C(_00484_),
    .D_N(net47),
    .X(_05121_));
 sky130_fd_sc_hd__a22o_1 _06024_ (.A1(net4),
    .A2(net46),
    .B1(net47),
    .B2(net3),
    .X(_05122_));
 sky130_fd_sc_hd__nand4_2 _06025_ (.A(_05121_),
    .B(net2),
    .C(net117),
    .D(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__a22o_1 _06026_ (.A1(net2),
    .A2(net117),
    .B1(_05121_),
    .B2(_05122_),
    .X(_05124_));
 sky130_fd_sc_hd__nand2_1 _06027_ (.A(_05123_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__and4_1 _06028_ (.A(net5),
    .B(net6),
    .C(net43),
    .D(net42),
    .X(_05126_));
 sky130_fd_sc_hd__o22a_1 _06029_ (.A1(_00154_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00187_),
    .X(_05127_));
 sky130_fd_sc_hd__a22o_1 _06030_ (.A1(net5),
    .A2(net43),
    .B1(net42),
    .B2(net6),
    .X(_05128_));
 sky130_fd_sc_hd__and4b_1 _06031_ (.A_N(_05126_),
    .B(_05128_),
    .C(net4),
    .D(net45),
    .X(_05129_));
 sky130_fd_sc_hd__a31o_1 _06032_ (.A1(_05128_),
    .A2(net45),
    .A3(net4),
    .B1(_05126_),
    .X(_05130_));
 sky130_fd_sc_hd__a22o_1 _06033_ (.A1(net5),
    .A2(net45),
    .B1(_05040_),
    .B2(_05041_),
    .X(_05131_));
 sky130_fd_sc_hd__and3_1 _06034_ (.A(_05042_),
    .B(_05130_),
    .C(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__a21oi_1 _06035_ (.A1(_05042_),
    .A2(_05131_),
    .B1(_05130_),
    .Y(_05133_));
 sky130_fd_sc_hd__nor2_1 _06036_ (.A(_05132_),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__xor2_1 _06037_ (.A(_05125_),
    .B(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__or2_1 _06038_ (.A(_05120_),
    .B(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__o21ai_1 _06039_ (.A1(_05120_),
    .A2(_05135_),
    .B1(_05119_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_1 _06040_ (.A(net14),
    .B(net64),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _06041_ (.A(net14),
    .B(net34),
    .Y(_05139_));
 sky130_fd_sc_hd__a22o_1 _06042_ (.A1(net15),
    .A2(net64),
    .B1(net34),
    .B2(net14),
    .X(_05140_));
 sky130_fd_sc_hd__nand3_1 _06043_ (.A(_05139_),
    .B(net64),
    .C(net15),
    .Y(_05141_));
 sky130_fd_sc_hd__nand3_1 _06044_ (.A(_05056_),
    .B(net34),
    .C(net14),
    .Y(_05142_));
 sky130_fd_sc_hd__o2111ai_4 _06045_ (.A1(_04985_),
    .A2(_05138_),
    .B1(net13),
    .C1(net35),
    .D1(_05140_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21ai_1 _06046_ (.A1(_04985_),
    .A2(_05138_),
    .B1(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__o2bb2a_1 _06047_ (.A1_N(_05057_),
    .A2_N(_05058_),
    .B1(_00242_),
    .B2(_00407_),
    .X(_05145_));
 sky130_fd_sc_hd__a22o_1 _06048_ (.A1(net14),
    .A2(net35),
    .B1(_05057_),
    .B2(_05058_),
    .X(_05146_));
 sky130_fd_sc_hd__nand3_1 _06049_ (.A(_05060_),
    .B(_05144_),
    .C(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__a21o_1 _06050_ (.A1(_05060_),
    .A2(_05146_),
    .B1(_05144_),
    .X(_05148_));
 sky130_fd_sc_hd__o21ai_1 _06051_ (.A1(_05059_),
    .A2(_05145_),
    .B1(_05144_),
    .Y(_05149_));
 sky130_fd_sc_hd__nand3b_1 _06052_ (.A_N(_05144_),
    .B(_05146_),
    .C(_05060_),
    .Y(_05150_));
 sky130_fd_sc_hd__o2bb2a_1 _06053_ (.A1_N(net10),
    .A2_N(net38),
    .B1(_05017_),
    .B2(_05018_),
    .X(_05151_));
 sky130_fd_sc_hd__nor2_1 _06054_ (.A(_05020_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand3_1 _06055_ (.A(_05147_),
    .B(_05148_),
    .C(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand3_1 _06056_ (.A(_05061_),
    .B(_05062_),
    .C(_05064_),
    .Y(_05154_));
 sky130_fd_sc_hd__a21o_1 _06057_ (.A1(_05061_),
    .A2(_05062_),
    .B1(_05064_),
    .X(_05155_));
 sky130_fd_sc_hd__nand2_1 _06058_ (.A(_05154_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__a21o_1 _06059_ (.A1(_05147_),
    .A2(_05153_),
    .B1(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__nand2_1 _06060_ (.A(_05033_),
    .B(_05050_),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_1 _06061_ (.A(_05051_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__xnor2_2 _06062_ (.A(_05157_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a21o_1 _06063_ (.A1(_05119_),
    .A2(_05136_),
    .B1(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__xnor2_2 _06064_ (.A(_05137_),
    .B(_05160_),
    .Y(_05162_));
 sky130_fd_sc_hd__inv_2 _06065_ (.A(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__or2_1 _06066_ (.A(_05053_),
    .B(_05065_),
    .X(_05164_));
 sky130_fd_sc_hd__nand2_2 _06067_ (.A(_05066_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__nor2_1 _06068_ (.A(_05163_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _06069_ (.A(_05016_),
    .B(_05073_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_1 _06070_ (.A(_05074_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nor2_1 _06071_ (.A(_05034_),
    .B(_05037_),
    .Y(_05169_));
 sky130_fd_sc_hd__a31o_1 _06072_ (.A1(_04974_),
    .A2(_05043_),
    .A3(_05044_),
    .B1(_05048_),
    .X(_05170_));
 sky130_fd_sc_hd__o21a_1 _06073_ (.A1(_05157_),
    .A2(_05159_),
    .B1(_05161_),
    .X(_05171_));
 sky130_fd_sc_hd__inv_2 _06074_ (.A(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _06075_ (.A(_05170_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a311o_1 _06076_ (.A1(_04974_),
    .A2(_05043_),
    .A3(_05044_),
    .B1(_05048_),
    .C1(_05172_),
    .X(_05174_));
 sky130_fd_sc_hd__nand2_1 _06077_ (.A(_05173_),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__xor2_1 _06078_ (.A(_05169_),
    .B(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__xnor2_1 _06079_ (.A(_05166_),
    .B(_05168_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2_1 _06080_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__o31ai_2 _06081_ (.A1(_05163_),
    .A2(_05165_),
    .A3(_05168_),
    .B1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _06082_ (.A(_05085_),
    .B(_05086_),
    .Y(_05180_));
 sky130_fd_sc_hd__xnor2_1 _06083_ (.A(_05085_),
    .B(_05086_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21ai_1 _06084_ (.A1(_05169_),
    .A2(_05175_),
    .B1(_05173_),
    .Y(_05182_));
 sky130_fd_sc_hd__xor2_1 _06085_ (.A(_05179_),
    .B(_05181_),
    .X(_05183_));
 sky130_fd_sc_hd__and2b_1 _06086_ (.A_N(_05183_),
    .B(_05182_),
    .X(_05184_));
 sky130_fd_sc_hd__a31o_1 _06087_ (.A1(_05087_),
    .A2(_05179_),
    .A3(_05180_),
    .B1(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__and2_1 _06088_ (.A(_05185_),
    .B(_05098_),
    .X(_05186_));
 sky130_fd_sc_hd__xnor2_1 _06089_ (.A(_05176_),
    .B(_05177_),
    .Y(_05187_));
 sky130_fd_sc_hd__xor2_1 _06090_ (.A(_05162_),
    .B(_05165_),
    .X(_05188_));
 sky130_fd_sc_hd__nand3_1 _06091_ (.A(_05156_),
    .B(_05153_),
    .C(_05147_),
    .Y(_05189_));
 sky130_fd_sc_hd__nand2_1 _06092_ (.A(_05157_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__and4_2 _06093_ (.A(net9),
    .B(net10),
    .C(net37),
    .D(net36),
    .X(_05191_));
 sky130_fd_sc_hd__o2bb2a_1 _06094_ (.A1_N(net9),
    .A2_N(net37),
    .B1(_00429_),
    .B2(_00231_),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _06095_ (.A1(net9),
    .A2(net37),
    .B1(net36),
    .B2(net10),
    .X(_05193_));
 sky130_fd_sc_hd__and4b_1 _06096_ (.A_N(_05191_),
    .B(_05193_),
    .C(net8),
    .D(net38),
    .X(_05194_));
 sky130_fd_sc_hd__a31oi_1 _06097_ (.A1(_05193_),
    .A2(net38),
    .A3(net8),
    .B1(_05191_),
    .Y(_05195_));
 sky130_fd_sc_hd__o22a_1 _06098_ (.A1(_00187_),
    .A2(_00451_),
    .B1(_05108_),
    .B2(_05109_),
    .X(_05196_));
 sky130_fd_sc_hd__nor2_1 _06099_ (.A(_05111_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__o21ai_4 _06100_ (.A1(_05191_),
    .A2(_05194_),
    .B1(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_1 _06101_ (.A(net6),
    .B(net39),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_1 _06102_ (.A(net6),
    .B(net40),
    .Y(_05200_));
 sky130_fd_sc_hd__a22o_1 _06103_ (.A1(net7),
    .A2(net39),
    .B1(net40),
    .B2(net6),
    .X(_05201_));
 sky130_fd_sc_hd__nand3_1 _06104_ (.A(_05200_),
    .B(net39),
    .C(net7),
    .Y(_05202_));
 sky130_fd_sc_hd__nand3_1 _06105_ (.A(_05106_),
    .B(net40),
    .C(net6),
    .Y(_05203_));
 sky130_fd_sc_hd__o2111ai_4 _06106_ (.A1(_05107_),
    .A2(_05199_),
    .B1(net5),
    .C1(net41),
    .D1(_05201_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21ai_2 _06107_ (.A1(_05106_),
    .A2(_05200_),
    .B1(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__o21ai_2 _06108_ (.A1(_05111_),
    .A2(_05196_),
    .B1(_05195_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand3_4 _06109_ (.A(_05198_),
    .B(_05205_),
    .C(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21oi_1 _06110_ (.A1(_05105_),
    .A2(_05113_),
    .B1(_05112_),
    .Y(_05208_));
 sky130_fd_sc_hd__a211o_1 _06111_ (.A1(_05198_),
    .A2(_05207_),
    .B1(_05208_),
    .C1(_05114_),
    .X(_05209_));
 sky130_fd_sc_hd__a22oi_1 _06112_ (.A1(net3),
    .A2(net46),
    .B1(net47),
    .B2(net2),
    .Y(_05210_));
 sky130_fd_sc_hd__and4_1 _06113_ (.A(net3),
    .B(net2),
    .C(net46),
    .D(net47),
    .X(_05211_));
 sky130_fd_sc_hd__o22a_1 _06114_ (.A1(_05210_),
    .A2(_05211_),
    .B1(_00110_),
    .B2(_00781_),
    .X(_05212_));
 sky130_fd_sc_hd__nor4_1 _06115_ (.A(_05210_),
    .B(_00110_),
    .C(_00781_),
    .D(_05211_),
    .Y(_05213_));
 sky130_fd_sc_hd__nand4_2 _06116_ (.A(net5),
    .B(net4),
    .C(net43),
    .D(net42),
    .Y(_05214_));
 sky130_fd_sc_hd__a22o_1 _06117_ (.A1(net4),
    .A2(net43),
    .B1(net42),
    .B2(net5),
    .X(_05215_));
 sky130_fd_sc_hd__and4_1 _06118_ (.A(_05215_),
    .B(net45),
    .C(net3),
    .D(_05214_),
    .X(_05216_));
 sky130_fd_sc_hd__nand4_1 _06119_ (.A(_05215_),
    .B(net45),
    .C(net3),
    .D(_05214_),
    .Y(_05217_));
 sky130_fd_sc_hd__o2bb2a_1 _06120_ (.A1_N(net4),
    .A2_N(net45),
    .B1(_05126_),
    .B2(_05127_),
    .X(_05218_));
 sky130_fd_sc_hd__o211ai_1 _06121_ (.A1(_05129_),
    .A2(_05218_),
    .B1(_05217_),
    .C1(_05214_),
    .Y(_05219_));
 sky130_fd_sc_hd__a211o_1 _06122_ (.A1(_05214_),
    .A2(_05217_),
    .B1(_05218_),
    .C1(_05129_),
    .X(_05220_));
 sky130_fd_sc_hd__a2bb2o_1 _06123_ (.A1_N(_05212_),
    .A2_N(_05213_),
    .B1(_05219_),
    .B2(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__or4bb_2 _06124_ (.A(_05212_),
    .B(_05213_),
    .C_N(_05219_),
    .D_N(_05220_),
    .X(_05222_));
 sky130_fd_sc_hd__o211ai_2 _06125_ (.A1(_05114_),
    .A2(_05208_),
    .B1(_05207_),
    .C1(_05198_),
    .Y(_05223_));
 sky130_fd_sc_hd__nand4_1 _06126_ (.A(_05209_),
    .B(_05221_),
    .C(_05222_),
    .D(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_1 _06127_ (.A(_05209_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__nand2_1 _06128_ (.A(_05120_),
    .B(_05135_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _06129_ (.A(_05136_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nor2_2 _06130_ (.A(_00264_),
    .B(_00374_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand2_2 _06131_ (.A(net15),
    .B(net62),
    .Y(_05229_));
 sky130_fd_sc_hd__or4_1 _06132_ (.A(_00264_),
    .B(_00374_),
    .C(_00396_),
    .D(_00869_),
    .X(_05230_));
 sky130_fd_sc_hd__o211ai_1 _06133_ (.A1(_05020_),
    .A2(_05151_),
    .B1(_05150_),
    .C1(_05149_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _06134_ (.A(_05153_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_1 _06135_ (.A(_05230_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__inv_2 _06136_ (.A(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(net13),
    .B(net64),
    .Y(_05235_));
 sky130_fd_sc_hd__nand4_1 _06138_ (.A(net14),
    .B(net13),
    .C(net64),
    .D(net34),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _06139_ (.A(net11),
    .B(net35),
    .Y(_05237_));
 sky130_fd_sc_hd__a22oi_1 _06140_ (.A1(net14),
    .A2(net64),
    .B1(net34),
    .B2(net13),
    .Y(_05238_));
 sky130_fd_sc_hd__a22o_1 _06141_ (.A1(net14),
    .A2(net64),
    .B1(net34),
    .B2(net13),
    .X(_05239_));
 sky130_fd_sc_hd__o2111ai_2 _06142_ (.A1(_05139_),
    .A2(_05235_),
    .B1(net11),
    .C1(net35),
    .D1(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ai_2 _06143_ (.A1(_05237_),
    .A2(_05238_),
    .B1(_05236_),
    .Y(_05241_));
 sky130_fd_sc_hd__o211ai_2 _06144_ (.A1(_00253_),
    .A2(_00407_),
    .B1(_05141_),
    .C1(_05142_),
    .Y(_05242_));
 sky130_fd_sc_hd__and3_1 _06145_ (.A(_05143_),
    .B(_05241_),
    .C(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__nand3_1 _06146_ (.A(_05143_),
    .B(_05241_),
    .C(_05242_),
    .Y(_05244_));
 sky130_fd_sc_hd__a2bb2o_1 _06147_ (.A1_N(_05099_),
    .A2_N(_05100_),
    .B1(net9),
    .B2(net38),
    .X(_05245_));
 sky130_fd_sc_hd__a21oi_1 _06148_ (.A1(_05143_),
    .A2(_05242_),
    .B1(_05241_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21o_1 _06149_ (.A1(_05143_),
    .A2(_05242_),
    .B1(_05241_),
    .X(_05247_));
 sky130_fd_sc_hd__nand4_1 _06150_ (.A(_05102_),
    .B(_05244_),
    .C(_05245_),
    .D(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__a31o_1 _06151_ (.A1(_05102_),
    .A2(_05245_),
    .A3(_05247_),
    .B1(_05243_),
    .X(_05249_));
 sky130_fd_sc_hd__a32o_1 _06152_ (.A1(net63),
    .A2(_05228_),
    .A3(net116),
    .B1(_05153_),
    .B2(_05231_),
    .X(_05250_));
 sky130_fd_sc_hd__nand3_1 _06153_ (.A(_05234_),
    .B(_05249_),
    .C(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__a21oi_1 _06154_ (.A1(_05234_),
    .A2(_05251_),
    .B1(_05227_),
    .Y(_05252_));
 sky130_fd_sc_hd__o211ai_1 _06155_ (.A1(_05230_),
    .A2(_05232_),
    .B1(_05251_),
    .C1(_05227_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2b_1 _06156_ (.A_N(_05252_),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__xor2_1 _06157_ (.A(_05225_),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__or2_1 _06158_ (.A(_05190_),
    .B(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__xor2_1 _06159_ (.A(_05188_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__a31o_1 _06160_ (.A1(_05134_),
    .A2(_05124_),
    .A3(_05123_),
    .B1(_05132_),
    .X(_05258_));
 sky130_fd_sc_hd__a21o_1 _06161_ (.A1(_05225_),
    .A2(_05253_),
    .B1(_05252_),
    .X(_05259_));
 sky130_fd_sc_hd__xnor2_1 _06162_ (.A(_05258_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__a21oi_1 _06163_ (.A1(_05121_),
    .A2(_05123_),
    .B1(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__and3_1 _06164_ (.A(_05121_),
    .B(_05123_),
    .C(_05260_),
    .X(_05262_));
 sky130_fd_sc_hd__nor2_1 _06165_ (.A(_05261_),
    .B(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand2_1 _06166_ (.A(_05257_),
    .B(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__o31a_1 _06167_ (.A1(_05188_),
    .A2(_05190_),
    .A3(_05255_),
    .B1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__or2_1 _06168_ (.A(_05265_),
    .B(_05187_),
    .X(_05266_));
 sky130_fd_sc_hd__a21oi_1 _06169_ (.A1(_05258_),
    .A2(_05259_),
    .B1(_05261_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _06170_ (.A(_05187_),
    .B(_05265_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _06171_ (.A(_05266_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21a_1 _06172_ (.A1(_05267_),
    .A2(_05269_),
    .B1(_05266_),
    .X(_05270_));
 sky130_fd_sc_hd__xor2_1 _06173_ (.A(_05182_),
    .B(_05183_),
    .X(_05271_));
 sky130_fd_sc_hd__nor2_1 _06174_ (.A(_05270_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__and2_1 _06175_ (.A(_05271_),
    .B(_05270_),
    .X(_05273_));
 sky130_fd_sc_hd__nor2_2 _06176_ (.A(_05272_),
    .B(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__a311o_1 _06177_ (.A1(net118),
    .A2(_00847_),
    .A3(_00000_),
    .B1(_00396_),
    .C1(_05228_),
    .X(_05275_));
 sky130_fd_sc_hd__nand2_1 _06178_ (.A(net11),
    .B(net34),
    .Y(_05276_));
 sky130_fd_sc_hd__nand4_1 _06179_ (.A(net11),
    .B(net13),
    .C(net64),
    .D(net34),
    .Y(_05277_));
 sky130_fd_sc_hd__a22o_1 _06180_ (.A1(net13),
    .A2(net64),
    .B1(net34),
    .B2(net11),
    .X(_05278_));
 sky130_fd_sc_hd__nand3_1 _06181_ (.A(_05276_),
    .B(net64),
    .C(net13),
    .Y(_05279_));
 sky130_fd_sc_hd__nand3_1 _06182_ (.A(_05235_),
    .B(net34),
    .C(net11),
    .Y(_05280_));
 sky130_fd_sc_hd__nand4_2 _06183_ (.A(_05278_),
    .B(net35),
    .C(net10),
    .D(_05277_),
    .Y(_05281_));
 sky130_fd_sc_hd__o21ai_1 _06184_ (.A1(_05235_),
    .A2(_05276_),
    .B1(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__a22o_1 _06185_ (.A1(net11),
    .A2(net35),
    .B1(_05236_),
    .B2(_05239_),
    .X(_05283_));
 sky130_fd_sc_hd__nand3_2 _06186_ (.A(_05240_),
    .B(_05282_),
    .C(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__a21o_1 _06187_ (.A1(_05240_),
    .A2(_05283_),
    .B1(_05282_),
    .X(_05285_));
 sky130_fd_sc_hd__o2bb2a_1 _06188_ (.A1_N(net8),
    .A2_N(net38),
    .B1(_05191_),
    .B2(_05192_),
    .X(_05286_));
 sky130_fd_sc_hd__a2bb2o_1 _06189_ (.A1_N(_05191_),
    .A2_N(_05192_),
    .B1(net8),
    .B2(net38),
    .X(_05287_));
 sky130_fd_sc_hd__nand4b_2 _06190_ (.A_N(_05194_),
    .B(_05284_),
    .C(_05285_),
    .D(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__a22oi_2 _06191_ (.A1(net15),
    .A2(net63),
    .B1(net116),
    .B2(net62),
    .Y(_05289_));
 sky130_fd_sc_hd__a31oi_4 _06192_ (.A1(net63),
    .A2(net116),
    .A3(_05228_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand4_2 _06193_ (.A(net116),
    .B(net61),
    .C(net62),
    .D(net15),
    .Y(_05291_));
 sky130_fd_sc_hd__nand2_1 _06194_ (.A(net14),
    .B(net63),
    .Y(_05292_));
 sky130_fd_sc_hd__a21oi_1 _06195_ (.A1(net116),
    .A2(net61),
    .B1(_05228_),
    .Y(_05293_));
 sky130_fd_sc_hd__o2bb2ai_1 _06196_ (.A1_N(net61),
    .A2_N(net116),
    .B1(_00264_),
    .B2(_00374_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand4_2 _06197_ (.A(_05294_),
    .B(net63),
    .C(net14),
    .D(_05291_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_2 _06198_ (.A1(_05292_),
    .A2(_05293_),
    .B1(_05291_),
    .Y(_05296_));
 sky130_fd_sc_hd__o2bb2ai_1 _06199_ (.A1_N(_05102_),
    .A2_N(_05245_),
    .B1(_05246_),
    .B2(_05243_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand4_2 _06200_ (.A(_05248_),
    .B(_05297_),
    .C(_05290_),
    .D(_05296_),
    .Y(_05298_));
 sky130_fd_sc_hd__a22o_1 _06201_ (.A1(_05290_),
    .A2(_05296_),
    .B1(_05297_),
    .B2(_05248_),
    .X(_05299_));
 sky130_fd_sc_hd__nand2_1 _06202_ (.A(_05298_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__a21o_1 _06203_ (.A1(_05284_),
    .A2(_05288_),
    .B1(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__nand3_1 _06204_ (.A(_05284_),
    .B(_05288_),
    .C(_05300_),
    .Y(_05302_));
 sky130_fd_sc_hd__and2_1 _06205_ (.A(_05301_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__and4_1 _06206_ (.A(net116),
    .B(_05303_),
    .C(_05229_),
    .D(net63),
    .X(_05304_));
 sky130_fd_sc_hd__a21o_1 _06207_ (.A1(_05234_),
    .A2(_05250_),
    .B1(_05249_),
    .X(_05305_));
 sky130_fd_sc_hd__nand2_1 _06208_ (.A(_05251_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__or4bb_1 _06209_ (.A(_05275_),
    .B(_05306_),
    .C_N(_05302_),
    .D_N(_05301_),
    .X(_05307_));
 sky130_fd_sc_hd__nand4_2 _06210_ (.A(net9),
    .B(net8),
    .C(net37),
    .D(net36),
    .Y(_05308_));
 sky130_fd_sc_hd__a22oi_1 _06211_ (.A1(net8),
    .A2(net37),
    .B1(net36),
    .B2(net9),
    .Y(_05309_));
 sky130_fd_sc_hd__a22o_1 _06212_ (.A1(net8),
    .A2(net37),
    .B1(net36),
    .B2(net9),
    .X(_05310_));
 sky130_fd_sc_hd__nand2_1 _06213_ (.A(net7),
    .B(net38),
    .Y(_05311_));
 sky130_fd_sc_hd__and4_1 _06214_ (.A(_05310_),
    .B(net38),
    .C(net7),
    .D(_05308_),
    .X(_05312_));
 sky130_fd_sc_hd__or3b_2 _06215_ (.A(_05311_),
    .B(_05309_),
    .C_N(_05308_),
    .X(_05313_));
 sky130_fd_sc_hd__o21ai_1 _06216_ (.A1(_05311_),
    .A2(_05309_),
    .B1(_05308_),
    .Y(_05314_));
 sky130_fd_sc_hd__o211ai_2 _06217_ (.A1(_00154_),
    .A2(_00451_),
    .B1(_05202_),
    .C1(_05203_),
    .Y(_05315_));
 sky130_fd_sc_hd__and3_1 _06218_ (.A(_05204_),
    .B(_05314_),
    .C(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__nand3_1 _06219_ (.A(_05204_),
    .B(_05314_),
    .C(_05315_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand2_2 _06220_ (.A(net5),
    .B(net40),
    .Y(_05318_));
 sky130_fd_sc_hd__nand4_2 _06221_ (.A(net5),
    .B(net6),
    .C(net39),
    .D(net40),
    .Y(_05319_));
 sky130_fd_sc_hd__a22o_1 _06222_ (.A1(net6),
    .A2(net39),
    .B1(net40),
    .B2(net5),
    .X(_05320_));
 sky130_fd_sc_hd__nand4_2 _06223_ (.A(_05320_),
    .B(net41),
    .C(net4),
    .D(_05319_),
    .Y(_05321_));
 sky130_fd_sc_hd__o21ai_1 _06224_ (.A1(_05199_),
    .A2(_05318_),
    .B1(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__a21o_1 _06225_ (.A1(_05204_),
    .A2(_05315_),
    .B1(_05314_),
    .X(_05323_));
 sky130_fd_sc_hd__and3_1 _06226_ (.A(_05317_),
    .B(_05322_),
    .C(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__a21o_1 _06227_ (.A1(_05198_),
    .A2(_05206_),
    .B1(_05205_),
    .X(_05325_));
 sky130_fd_sc_hd__o211ai_4 _06228_ (.A1(_05316_),
    .A2(_05324_),
    .B1(_05325_),
    .C1(_05207_),
    .Y(_05326_));
 sky130_fd_sc_hd__a22o_1 _06229_ (.A1(net2),
    .A2(net46),
    .B1(net47),
    .B2(net32),
    .X(_05327_));
 sky130_fd_sc_hd__or4b_2 _06230_ (.A(_00110_),
    .B(_00143_),
    .C(_00484_),
    .D_N(net47),
    .X(_05328_));
 sky130_fd_sc_hd__a22o_1 _06231_ (.A1(net117),
    .A2(net31),
    .B1(_05328_),
    .B2(_05327_),
    .X(_05329_));
 sky130_fd_sc_hd__nand4_2 _06232_ (.A(net117),
    .B(_05327_),
    .C(_05328_),
    .D(net31),
    .Y(_05330_));
 sky130_fd_sc_hd__nand4_4 _06233_ (.A(net3),
    .B(net4),
    .C(net43),
    .D(net42),
    .Y(_05331_));
 sky130_fd_sc_hd__a22o_1 _06234_ (.A1(net3),
    .A2(net43),
    .B1(net42),
    .B2(net4),
    .X(_05332_));
 sky130_fd_sc_hd__and4_1 _06235_ (.A(_05332_),
    .B(net45),
    .C(net2),
    .D(_05331_),
    .X(_05333_));
 sky130_fd_sc_hd__nand4_1 _06236_ (.A(_05332_),
    .B(net45),
    .C(net2),
    .D(_05331_),
    .Y(_05334_));
 sky130_fd_sc_hd__a22oi_2 _06237_ (.A1(net3),
    .A2(net45),
    .B1(_05214_),
    .B2(_05215_),
    .Y(_05335_));
 sky130_fd_sc_hd__o211ai_2 _06238_ (.A1(_05216_),
    .A2(_05335_),
    .B1(_05334_),
    .C1(_05331_),
    .Y(_05336_));
 sky130_fd_sc_hd__a211o_1 _06239_ (.A1(_05331_),
    .A2(_05334_),
    .B1(_05335_),
    .C1(_05216_),
    .X(_05337_));
 sky130_fd_sc_hd__a22o_1 _06240_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05336_),
    .B2(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__nand4_2 _06241_ (.A(_05329_),
    .B(_05330_),
    .C(_05336_),
    .D(_05337_),
    .Y(_05340_));
 sky130_fd_sc_hd__a221o_1 _06242_ (.A1(_05322_),
    .A2(_05323_),
    .B1(_05325_),
    .B2(_05207_),
    .C1(_05316_),
    .X(_05341_));
 sky130_fd_sc_hd__nand4_2 _06243_ (.A(_05326_),
    .B(_05338_),
    .C(_05340_),
    .D(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__nand2_1 _06244_ (.A(_05326_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__a22oi_1 _06245_ (.A1(_05221_),
    .A2(_05222_),
    .B1(_05223_),
    .B2(_05209_),
    .Y(_05344_));
 sky130_fd_sc_hd__a41o_1 _06246_ (.A1(_05209_),
    .A2(_05221_),
    .A3(_05222_),
    .A4(_05223_),
    .B1(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__a21o_1 _06247_ (.A1(_05298_),
    .A2(_05301_),
    .B1(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__nand3_1 _06248_ (.A(_05298_),
    .B(_05301_),
    .C(_05345_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__a21o_1 _06250_ (.A1(_05326_),
    .A2(_05342_),
    .B1(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__xnor2_1 _06251_ (.A(_05343_),
    .B(_05348_),
    .Y(_00001_));
 sky130_fd_sc_hd__xor2_2 _06252_ (.A(_05304_),
    .B(_05306_),
    .X(_00002_));
 sky130_fd_sc_hd__inv_2 _06253_ (.A(_00002_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_1 _06254_ (.A(_00001_),
    .B(_00003_),
    .Y(_00004_));
 sky130_fd_sc_hd__nand2_1 _06255_ (.A(_05190_),
    .B(_05255_),
    .Y(_00005_));
 sky130_fd_sc_hd__nand2_1 _06256_ (.A(_05256_),
    .B(_00005_),
    .Y(_00006_));
 sky130_fd_sc_hd__a21o_1 _06257_ (.A1(_05307_),
    .A2(_00004_),
    .B1(_00006_),
    .X(_00007_));
 sky130_fd_sc_hd__nand3_1 _06258_ (.A(_05307_),
    .B(_00004_),
    .C(_00006_),
    .Y(_00008_));
 sky130_fd_sc_hd__nand2_1 _06259_ (.A(_00007_),
    .B(_00008_),
    .Y(_00009_));
 sky130_fd_sc_hd__a41o_1 _06260_ (.A1(net3),
    .A2(net2),
    .A3(net46),
    .A4(net47),
    .B1(_05213_),
    .X(_00010_));
 sky130_fd_sc_hd__nand2_1 _06261_ (.A(_05220_),
    .B(_05222_),
    .Y(_00012_));
 sky130_fd_sc_hd__nand2_1 _06262_ (.A(_05346_),
    .B(_05349_),
    .Y(_00013_));
 sky130_fd_sc_hd__a22oi_1 _06263_ (.A1(_05220_),
    .A2(_05222_),
    .B1(_05346_),
    .B2(_05349_),
    .Y(_00014_));
 sky130_fd_sc_hd__and4_1 _06264_ (.A(_05220_),
    .B(_05222_),
    .C(_05346_),
    .D(_05349_),
    .X(_00015_));
 sky130_fd_sc_hd__nor2_1 _06265_ (.A(_00014_),
    .B(_00015_),
    .Y(_00016_));
 sky130_fd_sc_hd__o21a_1 _06266_ (.A1(_05211_),
    .A2(_05213_),
    .B1(_00016_),
    .X(_00017_));
 sky130_fd_sc_hd__nor2_1 _06267_ (.A(_00010_),
    .B(_00016_),
    .Y(_00018_));
 sky130_fd_sc_hd__or2_1 _06268_ (.A(_00017_),
    .B(_00018_),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _06269_ (.A(_00009_),
    .B(_00019_),
    .X(_00020_));
 sky130_fd_sc_hd__xnor2_1 _06270_ (.A(_05257_),
    .B(_05263_),
    .Y(_00021_));
 sky130_fd_sc_hd__a21o_1 _06271_ (.A1(_00007_),
    .A2(_00020_),
    .B1(_00021_),
    .X(_00023_));
 sky130_fd_sc_hd__o211ai_1 _06272_ (.A1(_00009_),
    .A2(_00019_),
    .B1(_00021_),
    .C1(_00007_),
    .Y(_00024_));
 sky130_fd_sc_hd__and2_1 _06273_ (.A(_00023_),
    .B(_00024_),
    .X(_00025_));
 sky130_fd_sc_hd__o21ai_1 _06274_ (.A1(_00014_),
    .A2(_00017_),
    .B1(_00025_),
    .Y(_00026_));
 sky130_fd_sc_hd__nand2_1 _06275_ (.A(_00023_),
    .B(_00026_),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _06276_ (.A(_00027_),
    .Y(_00028_));
 sky130_fd_sc_hd__xor2_1 _06277_ (.A(_05267_),
    .B(_05269_),
    .X(_00029_));
 sky130_fd_sc_hd__inv_2 _06278_ (.A(_00029_),
    .Y(_00030_));
 sky130_fd_sc_hd__or2_1 _06279_ (.A(_00027_),
    .B(_00029_),
    .X(_00031_));
 sky130_fd_sc_hd__a21o_1 _06280_ (.A1(_00023_),
    .A2(_00026_),
    .B1(_00030_),
    .X(_00032_));
 sky130_fd_sc_hd__a221o_1 _06281_ (.A1(_00012_),
    .A2(_00013_),
    .B1(_00016_),
    .B2(_00010_),
    .C1(_00025_),
    .X(_00034_));
 sky130_fd_sc_hd__nand2_1 _06282_ (.A(_00026_),
    .B(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__nand2_1 _06283_ (.A(net10),
    .B(net64),
    .Y(_00036_));
 sky130_fd_sc_hd__and4_1 _06284_ (.A(net11),
    .B(net10),
    .C(net64),
    .D(net34),
    .X(_00037_));
 sky130_fd_sc_hd__nand2_1 _06285_ (.A(net9),
    .B(net35),
    .Y(_00038_));
 sky130_fd_sc_hd__a22oi_2 _06286_ (.A1(net11),
    .A2(net64),
    .B1(net34),
    .B2(net10),
    .Y(_00039_));
 sky130_fd_sc_hd__a22o_1 _06287_ (.A1(net11),
    .A2(net64),
    .B1(net34),
    .B2(net10),
    .X(_00040_));
 sky130_fd_sc_hd__o2111ai_2 _06288_ (.A1(_05276_),
    .A2(_00036_),
    .B1(net9),
    .C1(net35),
    .D1(_00040_),
    .Y(_00041_));
 sky130_fd_sc_hd__o22ai_2 _06289_ (.A1(_05276_),
    .A2(_00036_),
    .B1(_00038_),
    .B2(_00039_),
    .Y(_00042_));
 sky130_fd_sc_hd__o211ai_2 _06290_ (.A1(_00231_),
    .A2(_00407_),
    .B1(_05279_),
    .C1(_05280_),
    .Y(_00043_));
 sky130_fd_sc_hd__and3_1 _06291_ (.A(_05281_),
    .B(_00042_),
    .C(_00043_),
    .X(_00045_));
 sky130_fd_sc_hd__nand3_1 _06292_ (.A(_05281_),
    .B(_00042_),
    .C(_00043_),
    .Y(_00046_));
 sky130_fd_sc_hd__a22oi_1 _06293_ (.A1(net7),
    .A2(net38),
    .B1(_05308_),
    .B2(_05310_),
    .Y(_00047_));
 sky130_fd_sc_hd__a22o_1 _06294_ (.A1(net7),
    .A2(net38),
    .B1(_05308_),
    .B2(_05310_),
    .X(_00048_));
 sky130_fd_sc_hd__a21oi_1 _06295_ (.A1(_05281_),
    .A2(_00043_),
    .B1(_00042_),
    .Y(_00049_));
 sky130_fd_sc_hd__a21o_1 _06296_ (.A1(_05281_),
    .A2(_00043_),
    .B1(_00042_),
    .X(_00050_));
 sky130_fd_sc_hd__nand4_1 _06297_ (.A(_05313_),
    .B(_00046_),
    .C(_00048_),
    .D(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__a31o_1 _06298_ (.A1(_05313_),
    .A2(_00048_),
    .A3(_00050_),
    .B1(_00045_),
    .X(_00052_));
 sky130_fd_sc_hd__o2bb2ai_2 _06299_ (.A1_N(_05291_),
    .A2_N(_05294_),
    .B1(_00242_),
    .B2(_00396_),
    .Y(_00053_));
 sky130_fd_sc_hd__nand2_1 _06300_ (.A(_05295_),
    .B(_00053_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand2_1 _06301_ (.A(net14),
    .B(net61),
    .Y(_00056_));
 sky130_fd_sc_hd__and3_1 _06302_ (.A(net14),
    .B(net61),
    .C(_05228_),
    .X(_00057_));
 sky130_fd_sc_hd__nand4_1 _06303_ (.A(net14),
    .B(net15),
    .C(net62),
    .D(net61),
    .Y(_00058_));
 sky130_fd_sc_hd__a22o_2 _06304_ (.A1(net14),
    .A2(net62),
    .B1(net61),
    .B2(net15),
    .X(_00059_));
 sky130_fd_sc_hd__o2111a_2 _06305_ (.A1(_05229_),
    .A2(_00056_),
    .B1(net13),
    .C1(net63),
    .D1(_00059_),
    .X(_00060_));
 sky130_fd_sc_hd__o2111ai_4 _06306_ (.A1(_05229_),
    .A2(_00056_),
    .B1(net13),
    .C1(net63),
    .D1(_00059_),
    .Y(_00061_));
 sky130_fd_sc_hd__o31a_1 _06307_ (.A1(_00242_),
    .A2(_00385_),
    .A3(_05229_),
    .B1(_00061_),
    .X(_00062_));
 sky130_fd_sc_hd__o211ai_4 _06308_ (.A1(_00057_),
    .A2(_00060_),
    .B1(_05295_),
    .C1(_00053_),
    .Y(_00063_));
 sky130_fd_sc_hd__o2bb2ai_1 _06309_ (.A1_N(_05284_),
    .A2_N(_05285_),
    .B1(_05286_),
    .B2(_05194_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand3b_1 _06310_ (.A_N(_00063_),
    .B(_00064_),
    .C(_05288_),
    .Y(_00065_));
 sky130_fd_sc_hd__o2bb2ai_1 _06311_ (.A1_N(_05288_),
    .A2_N(_00064_),
    .B1(_00062_),
    .B2(_00054_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand3_1 _06312_ (.A(_00052_),
    .B(_00065_),
    .C(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__a21o_1 _06313_ (.A1(_00065_),
    .A2(_00067_),
    .B1(_00052_),
    .X(_00069_));
 sky130_fd_sc_hd__xor2_2 _06314_ (.A(_05290_),
    .B(_05296_),
    .X(_00070_));
 sky130_fd_sc_hd__nand3_1 _06315_ (.A(_00068_),
    .B(_00069_),
    .C(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__xnor2_1 _06316_ (.A(_05275_),
    .B(_05303_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand4_2 _06317_ (.A(net7),
    .B(net8),
    .C(net37),
    .D(net36),
    .Y(_00073_));
 sky130_fd_sc_hd__a22o_1 _06318_ (.A1(net7),
    .A2(net37),
    .B1(net36),
    .B2(net8),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _06319_ (.A(net6),
    .B(net38),
    .X(_00075_));
 sky130_fd_sc_hd__nand4_2 _06320_ (.A(_00074_),
    .B(net38),
    .C(net6),
    .D(_00073_),
    .Y(_00076_));
 sky130_fd_sc_hd__a21bo_1 _06321_ (.A1(_00074_),
    .A2(_00075_),
    .B1_N(_00073_),
    .X(_00078_));
 sky130_fd_sc_hd__o2bb2ai_1 _06322_ (.A1_N(_05319_),
    .A2_N(_05320_),
    .B1(_00165_),
    .B2(_00451_),
    .Y(_00079_));
 sky130_fd_sc_hd__nand3_1 _06323_ (.A(_05321_),
    .B(_00078_),
    .C(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_2 _06324_ (.A(net4),
    .B(net39),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(net4),
    .B(net40),
    .Y(_00082_));
 sky130_fd_sc_hd__nand4_1 _06326_ (.A(net5),
    .B(net4),
    .C(net39),
    .D(net40),
    .Y(_00083_));
 sky130_fd_sc_hd__a22o_1 _06327_ (.A1(net5),
    .A2(net39),
    .B1(net40),
    .B2(net4),
    .X(_00084_));
 sky130_fd_sc_hd__o2111ai_4 _06328_ (.A1(_05318_),
    .A2(_00081_),
    .B1(net3),
    .C1(net41),
    .D1(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__o21ai_1 _06329_ (.A1(_05318_),
    .A2(_00081_),
    .B1(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__a21o_1 _06330_ (.A1(_05321_),
    .A2(_00079_),
    .B1(_00078_),
    .X(_00087_));
 sky130_fd_sc_hd__nand3_1 _06331_ (.A(_00080_),
    .B(_00086_),
    .C(_00087_),
    .Y(_00089_));
 sky130_fd_sc_hd__a21boi_1 _06332_ (.A1(_00086_),
    .A2(_00087_),
    .B1_N(_00080_),
    .Y(_00090_));
 sky130_fd_sc_hd__a22o_1 _06333_ (.A1(_05319_),
    .A2(_05321_),
    .B1(_05323_),
    .B2(_05317_),
    .X(_00091_));
 sky130_fd_sc_hd__nand3b_1 _06334_ (.A_N(_05322_),
    .B(_05323_),
    .C(_05317_),
    .Y(_00092_));
 sky130_fd_sc_hd__a21oi_1 _06335_ (.A1(_00091_),
    .A2(_00092_),
    .B1(_00090_),
    .Y(_00093_));
 sky130_fd_sc_hd__a22o_1 _06336_ (.A1(net32),
    .A2(net46),
    .B1(net47),
    .B2(net31),
    .X(_00094_));
 sky130_fd_sc_hd__nand4_2 _06337_ (.A(net32),
    .B(net31),
    .C(net46),
    .D(net47),
    .Y(_00095_));
 sky130_fd_sc_hd__a22o_1 _06338_ (.A1(_00094_),
    .A2(_00095_),
    .B1(net117),
    .B2(net30),
    .X(_00096_));
 sky130_fd_sc_hd__nand4_2 _06339_ (.A(net117),
    .B(_00094_),
    .C(_00095_),
    .D(net30),
    .Y(_00097_));
 sky130_fd_sc_hd__nand4_4 _06340_ (.A(net3),
    .B(net2),
    .C(net43),
    .D(net42),
    .Y(_00098_));
 sky130_fd_sc_hd__a22o_1 _06341_ (.A1(net2),
    .A2(net43),
    .B1(net42),
    .B2(net3),
    .X(_00100_));
 sky130_fd_sc_hd__and4_1 _06342_ (.A(_00100_),
    .B(net45),
    .C(net32),
    .D(_00098_),
    .X(_00101_));
 sky130_fd_sc_hd__nand4_1 _06343_ (.A(_00100_),
    .B(net45),
    .C(net32),
    .D(_00098_),
    .Y(_00102_));
 sky130_fd_sc_hd__a22oi_2 _06344_ (.A1(net2),
    .A2(net45),
    .B1(_05331_),
    .B2(_05332_),
    .Y(_00103_));
 sky130_fd_sc_hd__o211ai_2 _06345_ (.A1(_05333_),
    .A2(_00103_),
    .B1(_00102_),
    .C1(_00098_),
    .Y(_00104_));
 sky130_fd_sc_hd__a211o_1 _06346_ (.A1(_00098_),
    .A2(_00102_),
    .B1(_00103_),
    .C1(_05333_),
    .X(_00105_));
 sky130_fd_sc_hd__a22o_1 _06347_ (.A1(_00096_),
    .A2(_00097_),
    .B1(_00104_),
    .B2(_00105_),
    .X(_00106_));
 sky130_fd_sc_hd__nand4_2 _06348_ (.A(_00096_),
    .B(_00097_),
    .C(_00104_),
    .D(_00105_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3_1 _06349_ (.A(_00090_),
    .B(_00091_),
    .C(_00092_),
    .X(_00108_));
 sky130_fd_sc_hd__nand4_1 _06350_ (.A(_00080_),
    .B(_00089_),
    .C(_00091_),
    .D(_00092_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand4b_1 _06351_ (.A_N(_00093_),
    .B(_00106_),
    .C(_00107_),
    .D(_00109_),
    .Y(_00111_));
 sky130_fd_sc_hd__a31o_1 _06352_ (.A1(_00106_),
    .A2(_00107_),
    .A3(_00109_),
    .B1(_00093_),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _06353_ (.A(_00065_),
    .B(_00068_),
    .Y(_00113_));
 sky130_fd_sc_hd__a22o_1 _06354_ (.A1(_05338_),
    .A2(_05340_),
    .B1(_05341_),
    .B2(_05326_),
    .X(_00114_));
 sky130_fd_sc_hd__nand3_1 _06355_ (.A(_05342_),
    .B(_00113_),
    .C(_00114_),
    .Y(_00115_));
 sky130_fd_sc_hd__a21o_1 _06356_ (.A1(_05342_),
    .A2(_00114_),
    .B1(_00113_),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _06357_ (.A(_00115_),
    .B(_00116_),
    .Y(_00117_));
 sky130_fd_sc_hd__xor2_1 _06358_ (.A(_00112_),
    .B(_00117_),
    .X(_00118_));
 sky130_fd_sc_hd__xor2_1 _06359_ (.A(_00071_),
    .B(_00072_),
    .X(_00119_));
 sky130_fd_sc_hd__nor2_1 _06360_ (.A(_00118_),
    .B(_00119_),
    .Y(_00120_));
 sky130_fd_sc_hd__a41o_1 _06361_ (.A1(_00068_),
    .A2(_00069_),
    .A3(_00070_),
    .A4(_00072_),
    .B1(_00120_),
    .X(_00122_));
 sky130_fd_sc_hd__xnor2_1 _06362_ (.A(_00001_),
    .B(_00002_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _06363_ (.A(_00123_),
    .B(_00122_),
    .Y(_00124_));
 sky130_fd_sc_hd__xnor2_1 _06364_ (.A(_00122_),
    .B(_00123_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _06365_ (.A(_05328_),
    .B(_05330_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _06366_ (.A(_05337_),
    .B(_05340_),
    .Y(_00127_));
 sky130_fd_sc_hd__a21bo_1 _06367_ (.A1(_00112_),
    .A2(_00116_),
    .B1_N(_00115_),
    .X(_00128_));
 sky130_fd_sc_hd__xor2_1 _06368_ (.A(_00127_),
    .B(_00128_),
    .X(_00129_));
 sky130_fd_sc_hd__xnor2_1 _06369_ (.A(_00126_),
    .B(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__o21a_1 _06370_ (.A1(_00125_),
    .A2(_00130_),
    .B1(_00124_),
    .X(_00131_));
 sky130_fd_sc_hd__nand2_1 _06371_ (.A(_00009_),
    .B(_00019_),
    .Y(_00133_));
 sky130_fd_sc_hd__nand2_1 _06372_ (.A(_00020_),
    .B(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__or2_1 _06373_ (.A(_00131_),
    .B(_00134_),
    .X(_00135_));
 sky130_fd_sc_hd__a22oi_2 _06374_ (.A1(_00127_),
    .A2(_00128_),
    .B1(_00129_),
    .B2(_00126_),
    .Y(_00136_));
 sky130_fd_sc_hd__xnor2_1 _06375_ (.A(_00131_),
    .B(_00134_),
    .Y(_00137_));
 sky130_fd_sc_hd__or2_1 _06376_ (.A(_00136_),
    .B(_00137_),
    .X(_00138_));
 sky130_fd_sc_hd__a21o_1 _06377_ (.A1(_00135_),
    .A2(_00138_),
    .B1(_00035_),
    .X(_00139_));
 sky130_fd_sc_hd__o211ai_2 _06378_ (.A1(_00131_),
    .A2(_00134_),
    .B1(_00138_),
    .C1(_00035_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand2_2 _06379_ (.A(_00139_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__a21bo_1 _06380_ (.A1(_05295_),
    .A2(_00053_),
    .B1_N(_00062_),
    .X(_00142_));
 sky130_fd_sc_hd__a21oi_4 _06381_ (.A1(net118),
    .A2(_00858_),
    .B1(_00352_),
    .Y(_00144_));
 sky130_fd_sc_hd__a31o_1 _06382_ (.A1(net118),
    .A2(_00847_),
    .A3(_00000_),
    .B1(_00352_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(net13),
    .B(net61),
    .Y(_00146_));
 sky130_fd_sc_hd__and4_1 _06384_ (.A(net14),
    .B(net13),
    .C(net62),
    .D(net61),
    .X(_00147_));
 sky130_fd_sc_hd__nand4_4 _06385_ (.A(net14),
    .B(net13),
    .C(net62),
    .D(net61),
    .Y(_00148_));
 sky130_fd_sc_hd__a22o_1 _06386_ (.A1(net13),
    .A2(net62),
    .B1(net61),
    .B2(net14),
    .X(_00149_));
 sky130_fd_sc_hd__and4_1 _06387_ (.A(_00149_),
    .B(net63),
    .C(net11),
    .D(_00148_),
    .X(_00150_));
 sky130_fd_sc_hd__nand4_2 _06388_ (.A(_00149_),
    .B(net63),
    .C(net11),
    .D(_00148_),
    .Y(_00151_));
 sky130_fd_sc_hd__o31a_1 _06389_ (.A1(_00242_),
    .A2(_00374_),
    .A3(_00146_),
    .B1(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__nor2_1 _06390_ (.A(_00264_),
    .B(_00363_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_2 _06391_ (.A(net15),
    .B(net59),
    .Y(_00155_));
 sky130_fd_sc_hd__nand4_2 _06392_ (.A(net116),
    .B(net59),
    .C(net60),
    .D(net15),
    .Y(_00156_));
 sky130_fd_sc_hd__a22oi_2 _06393_ (.A1(net13),
    .A2(net63),
    .B1(_00058_),
    .B2(_00059_),
    .Y(_00157_));
 sky130_fd_sc_hd__a22o_1 _06394_ (.A1(net13),
    .A2(net63),
    .B1(_00058_),
    .B2(_00059_),
    .X(_00158_));
 sky130_fd_sc_hd__nand4_4 _06395_ (.A(_00144_),
    .B(_00158_),
    .C(_00153_),
    .D(_00061_),
    .Y(_00159_));
 sky130_fd_sc_hd__o21ai_4 _06396_ (.A1(_00060_),
    .A2(_00157_),
    .B1(_00156_),
    .Y(_00160_));
 sky130_fd_sc_hd__o211ai_4 _06397_ (.A1(_00147_),
    .A2(_00150_),
    .B1(_00159_),
    .C1(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__a21bo_1 _06398_ (.A1(_00159_),
    .A2(_00160_),
    .B1_N(_00152_),
    .X(_00162_));
 sky130_fd_sc_hd__nand4_1 _06399_ (.A(_00148_),
    .B(_00151_),
    .C(_00159_),
    .D(_00160_),
    .Y(_00163_));
 sky130_fd_sc_hd__a22o_1 _06400_ (.A1(_00148_),
    .A2(_00151_),
    .B1(_00159_),
    .B2(_00160_),
    .X(_00164_));
 sky130_fd_sc_hd__nand2_1 _06401_ (.A(_00163_),
    .B(_00164_),
    .Y(_00166_));
 sky130_fd_sc_hd__a21o_1 _06402_ (.A1(_00163_),
    .A2(_00164_),
    .B1(_00145_),
    .X(_00167_));
 sky130_fd_sc_hd__nand4_1 _06403_ (.A(_00063_),
    .B(_00142_),
    .C(_00161_),
    .D(_00162_),
    .Y(_00168_));
 sky130_fd_sc_hd__a311o_1 _06404_ (.A1(_00000_),
    .A2(net118),
    .A3(_00847_),
    .B1(_00168_),
    .C1(_00352_),
    .X(_00169_));
 sky130_fd_sc_hd__a32o_1 _06405_ (.A1(_00144_),
    .A2(_00161_),
    .A3(_00162_),
    .B1(_00142_),
    .B2(_00063_),
    .X(_00170_));
 sky130_fd_sc_hd__nand2_1 _06406_ (.A(net9),
    .B(net64),
    .Y(_00171_));
 sky130_fd_sc_hd__and4_1 _06407_ (.A(net9),
    .B(net10),
    .C(net64),
    .D(net34),
    .X(_00172_));
 sky130_fd_sc_hd__a22oi_1 _06408_ (.A1(net10),
    .A2(net64),
    .B1(net34),
    .B2(net9),
    .Y(_00173_));
 sky130_fd_sc_hd__a22o_1 _06409_ (.A1(net10),
    .A2(net64),
    .B1(net34),
    .B2(net9),
    .X(_00174_));
 sky130_fd_sc_hd__nand4b_1 _06410_ (.A_N(_00172_),
    .B(_00174_),
    .C(net8),
    .D(net35),
    .Y(_00175_));
 sky130_fd_sc_hd__a31o_1 _06411_ (.A1(_00174_),
    .A2(net35),
    .A3(net8),
    .B1(_00172_),
    .X(_00177_));
 sky130_fd_sc_hd__o21ai_1 _06412_ (.A1(_00037_),
    .A2(_00039_),
    .B1(_00038_),
    .Y(_00178_));
 sky130_fd_sc_hd__and3_1 _06413_ (.A(_00041_),
    .B(_00177_),
    .C(_00178_),
    .X(_00179_));
 sky130_fd_sc_hd__nand3_1 _06414_ (.A(_00041_),
    .B(_00177_),
    .C(_00178_),
    .Y(_00180_));
 sky130_fd_sc_hd__a22o_1 _06415_ (.A1(net6),
    .A2(net38),
    .B1(_00073_),
    .B2(_00074_),
    .X(_00181_));
 sky130_fd_sc_hd__nand2_1 _06416_ (.A(_00076_),
    .B(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__a21o_1 _06417_ (.A1(_00041_),
    .A2(_00178_),
    .B1(_00177_),
    .X(_00183_));
 sky130_fd_sc_hd__and4_2 _06418_ (.A(_00076_),
    .B(_00180_),
    .C(_00181_),
    .D(_00183_),
    .X(_00184_));
 sky130_fd_sc_hd__a31o_1 _06419_ (.A1(_00076_),
    .A2(_00181_),
    .A3(_00183_),
    .B1(_00179_),
    .X(_00185_));
 sky130_fd_sc_hd__nand2_1 _06420_ (.A(_00159_),
    .B(_00161_),
    .Y(_00186_));
 sky130_fd_sc_hd__a22o_1 _06421_ (.A1(_05313_),
    .A2(_00048_),
    .B1(_00050_),
    .B2(_00046_),
    .X(_00188_));
 sky130_fd_sc_hd__o211ai_2 _06422_ (.A1(_00045_),
    .A2(_00049_),
    .B1(_00048_),
    .C1(_05313_),
    .Y(_00189_));
 sky130_fd_sc_hd__o211ai_2 _06423_ (.A1(_05312_),
    .A2(_00047_),
    .B1(_00050_),
    .C1(_00046_),
    .Y(_00190_));
 sky130_fd_sc_hd__a22oi_2 _06424_ (.A1(_00159_),
    .A2(_00161_),
    .B1(_00189_),
    .B2(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__a22o_1 _06425_ (.A1(_00159_),
    .A2(_00161_),
    .B1(_00189_),
    .B2(_00190_),
    .X(_00192_));
 sky130_fd_sc_hd__a21oi_1 _06426_ (.A1(_00051_),
    .A2(_00188_),
    .B1(_00186_),
    .Y(_00193_));
 sky130_fd_sc_hd__a21o_1 _06427_ (.A1(_00051_),
    .A2(_00188_),
    .B1(_00186_),
    .X(_00194_));
 sky130_fd_sc_hd__o211ai_4 _06428_ (.A1(_00179_),
    .A2(_00184_),
    .B1(_00192_),
    .C1(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__o21bai_2 _06429_ (.A1(_00191_),
    .A2(_00193_),
    .B1_N(_00185_),
    .Y(_00196_));
 sky130_fd_sc_hd__o2111a_2 _06430_ (.A1(_00145_),
    .A2(_00168_),
    .B1(_00170_),
    .C1(_00195_),
    .D1(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__a41oi_4 _06431_ (.A1(_00063_),
    .A2(_00142_),
    .A3(_00144_),
    .A4(_00166_),
    .B1(_00197_),
    .Y(_00199_));
 sky130_fd_sc_hd__a21o_1 _06432_ (.A1(_00068_),
    .A2(_00069_),
    .B1(_00070_),
    .X(_00200_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(_00071_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__xor2_1 _06434_ (.A(_00199_),
    .B(_00201_),
    .X(_00202_));
 sky130_fd_sc_hd__nand4_2 _06435_ (.A(net7),
    .B(net6),
    .C(net37),
    .D(net36),
    .Y(_00203_));
 sky130_fd_sc_hd__a22o_1 _06436_ (.A1(net6),
    .A2(net37),
    .B1(net36),
    .B2(net7),
    .X(_00204_));
 sky130_fd_sc_hd__nand4_2 _06437_ (.A(_00204_),
    .B(net38),
    .C(net5),
    .D(_00203_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(_00203_),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__a22o_1 _06439_ (.A1(net3),
    .A2(net41),
    .B1(_00083_),
    .B2(_00084_),
    .X(_00207_));
 sky130_fd_sc_hd__nand3_1 _06440_ (.A(_00085_),
    .B(_00206_),
    .C(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(net3),
    .B(net39),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _06442_ (.A(net3),
    .B(net40),
    .Y(_00211_));
 sky130_fd_sc_hd__a22o_1 _06443_ (.A1(net4),
    .A2(net39),
    .B1(net40),
    .B2(net3),
    .X(_00212_));
 sky130_fd_sc_hd__nand3_1 _06444_ (.A(_00211_),
    .B(net39),
    .C(net4),
    .Y(_00213_));
 sky130_fd_sc_hd__nand3_1 _06445_ (.A(_00081_),
    .B(net40),
    .C(net3),
    .Y(_00214_));
 sky130_fd_sc_hd__o2111ai_4 _06446_ (.A1(_00082_),
    .A2(_00210_),
    .B1(net2),
    .C1(net41),
    .D1(_00212_),
    .Y(_00215_));
 sky130_fd_sc_hd__o31a_1 _06447_ (.A1(_00165_),
    .A2(_00440_),
    .A3(_00211_),
    .B1(_00215_),
    .X(_00216_));
 sky130_fd_sc_hd__a21oi_1 _06448_ (.A1(_00085_),
    .A2(_00207_),
    .B1(_00206_),
    .Y(_00217_));
 sky130_fd_sc_hd__a21o_1 _06449_ (.A1(_00085_),
    .A2(_00207_),
    .B1(_00206_),
    .X(_00218_));
 sky130_fd_sc_hd__o21ai_1 _06450_ (.A1(_00216_),
    .A2(_00217_),
    .B1(_00208_),
    .Y(_00219_));
 sky130_fd_sc_hd__a21o_1 _06451_ (.A1(_00080_),
    .A2(_00087_),
    .B1(_00086_),
    .X(_00221_));
 sky130_fd_sc_hd__nand3_1 _06452_ (.A(_00089_),
    .B(_00219_),
    .C(_00221_),
    .Y(_00222_));
 sky130_fd_sc_hd__a21o_1 _06453_ (.A1(_00089_),
    .A2(_00221_),
    .B1(_00219_),
    .X(_00223_));
 sky130_fd_sc_hd__a22o_1 _06454_ (.A1(net31),
    .A2(net46),
    .B1(net47),
    .B2(net30),
    .X(_00224_));
 sky130_fd_sc_hd__nand4_2 _06455_ (.A(net30),
    .B(net31),
    .C(net46),
    .D(net47),
    .Y(_00225_));
 sky130_fd_sc_hd__a22o_1 _06456_ (.A1(_00224_),
    .A2(_00225_),
    .B1(net117),
    .B2(net29),
    .X(_00226_));
 sky130_fd_sc_hd__nand4_2 _06457_ (.A(net117),
    .B(_00224_),
    .C(_00225_),
    .D(net29),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _06458_ (.A(_00226_),
    .B(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand4_4 _06459_ (.A(net32),
    .B(net2),
    .C(net43),
    .D(net42),
    .Y(_00229_));
 sky130_fd_sc_hd__a22o_1 _06460_ (.A1(net32),
    .A2(net43),
    .B1(net42),
    .B2(net2),
    .X(_00230_));
 sky130_fd_sc_hd__nand4_4 _06461_ (.A(_00230_),
    .B(net45),
    .C(net31),
    .D(_00229_),
    .Y(_00232_));
 sky130_fd_sc_hd__a22oi_2 _06462_ (.A1(net32),
    .A2(net45),
    .B1(_00098_),
    .B2(_00100_),
    .Y(_00233_));
 sky130_fd_sc_hd__o211ai_2 _06463_ (.A1(_00101_),
    .A2(_00233_),
    .B1(_00232_),
    .C1(_00229_),
    .Y(_00234_));
 sky130_fd_sc_hd__a211o_1 _06464_ (.A1(_00229_),
    .A2(_00232_),
    .B1(_00233_),
    .C1(_00101_),
    .X(_00235_));
 sky130_fd_sc_hd__nand2_1 _06465_ (.A(_00234_),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__and4_1 _06466_ (.A(_00226_),
    .B(_00227_),
    .C(_00234_),
    .D(_00235_),
    .X(_00237_));
 sky130_fd_sc_hd__or2_1 _06467_ (.A(_00228_),
    .B(_00236_),
    .X(_00238_));
 sky130_fd_sc_hd__a22oi_1 _06468_ (.A1(_00226_),
    .A2(_00227_),
    .B1(_00234_),
    .B2(_00235_),
    .Y(_00239_));
 sky130_fd_sc_hd__a22o_1 _06469_ (.A1(_00226_),
    .A2(_00227_),
    .B1(_00234_),
    .B2(_00235_),
    .X(_00240_));
 sky130_fd_sc_hd__nand4_1 _06470_ (.A(_00222_),
    .B(_00223_),
    .C(_00238_),
    .D(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _06471_ (.A(_00222_),
    .B(_00241_),
    .Y(_00243_));
 sky130_fd_sc_hd__o2bb2ai_1 _06472_ (.A1_N(_00106_),
    .A2_N(_00107_),
    .B1(_00108_),
    .B2(_00093_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _06473_ (.A(_00111_),
    .B(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__a21oi_1 _06474_ (.A1(_00192_),
    .A2(_00195_),
    .B1(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__a221oi_1 _06475_ (.A1(_00185_),
    .A2(_00194_),
    .B1(_00244_),
    .B2(_00111_),
    .C1(_00191_),
    .Y(_00247_));
 sky130_fd_sc_hd__nor2_1 _06476_ (.A(_00246_),
    .B(_00247_),
    .Y(_00248_));
 sky130_fd_sc_hd__xor2_1 _06477_ (.A(_00243_),
    .B(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(_00202_),
    .B(_00249_),
    .Y(_00250_));
 sky130_fd_sc_hd__o21ai_1 _06479_ (.A1(_00199_),
    .A2(_00201_),
    .B1(_00250_),
    .Y(_00251_));
 sky130_fd_sc_hd__and2_1 _06480_ (.A(_00118_),
    .B(_00119_),
    .X(_00252_));
 sky130_fd_sc_hd__nor2_1 _06481_ (.A(_00120_),
    .B(_00252_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _06482_ (.A(_00095_),
    .B(_00097_),
    .Y(_00255_));
 sky130_fd_sc_hd__a21oi_1 _06483_ (.A1(_00248_),
    .A2(_00243_),
    .B1(_00246_),
    .Y(_00256_));
 sky130_fd_sc_hd__a21oi_1 _06484_ (.A1(_00105_),
    .A2(_00107_),
    .B1(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__and3_1 _06485_ (.A(_00256_),
    .B(_00107_),
    .C(_00105_),
    .X(_00258_));
 sky130_fd_sc_hd__nor2_1 _06486_ (.A(_00257_),
    .B(_00258_),
    .Y(_00259_));
 sky130_fd_sc_hd__xnor2_1 _06487_ (.A(_00255_),
    .B(_00259_),
    .Y(_00260_));
 sky130_fd_sc_hd__xor2_1 _06488_ (.A(_00251_),
    .B(_00254_),
    .X(_00261_));
 sky130_fd_sc_hd__and2b_1 _06489_ (.A_N(_00260_),
    .B(_00261_),
    .X(_00262_));
 sky130_fd_sc_hd__a21o_1 _06490_ (.A1(_00251_),
    .A2(_00254_),
    .B1(_00262_),
    .X(_00263_));
 sky130_fd_sc_hd__xnor2_1 _06491_ (.A(_00125_),
    .B(_00130_),
    .Y(_00265_));
 sky130_fd_sc_hd__and2b_1 _06492_ (.A_N(_00265_),
    .B(_00263_),
    .X(_00266_));
 sky130_fd_sc_hd__a21oi_1 _06493_ (.A1(_00259_),
    .A2(_00255_),
    .B1(_00257_),
    .Y(_00267_));
 sky130_fd_sc_hd__xor2_1 _06494_ (.A(_00263_),
    .B(_00265_),
    .X(_00268_));
 sky130_fd_sc_hd__o21bai_2 _06495_ (.A1(_00267_),
    .A2(_00268_),
    .B1_N(_00266_),
    .Y(_00269_));
 sky130_fd_sc_hd__xnor2_1 _06496_ (.A(_00136_),
    .B(_00137_),
    .Y(_00270_));
 sky130_fd_sc_hd__and2b_1 _06497_ (.A_N(_00270_),
    .B(_00269_),
    .X(_00271_));
 sky130_fd_sc_hd__a22o_1 _06498_ (.A1(net116),
    .A2(net60),
    .B1(_00162_),
    .B2(_00161_),
    .X(_00272_));
 sky130_fd_sc_hd__nand2_1 _06499_ (.A(net11),
    .B(net62),
    .Y(_00273_));
 sky130_fd_sc_hd__nand4_1 _06500_ (.A(net11),
    .B(net13),
    .C(net62),
    .D(net61),
    .Y(_00274_));
 sky130_fd_sc_hd__a22o_1 _06501_ (.A1(net11),
    .A2(net62),
    .B1(net61),
    .B2(net13),
    .X(_00276_));
 sky130_fd_sc_hd__nand3_1 _06502_ (.A(_00273_),
    .B(net61),
    .C(net13),
    .Y(_00277_));
 sky130_fd_sc_hd__nand3_1 _06503_ (.A(_00146_),
    .B(net62),
    .C(net11),
    .Y(_00278_));
 sky130_fd_sc_hd__nand4_2 _06504_ (.A(_00276_),
    .B(net63),
    .C(net10),
    .D(_00274_),
    .Y(_00279_));
 sky130_fd_sc_hd__o31a_2 _06505_ (.A1(_00220_),
    .A2(_00374_),
    .A3(_00146_),
    .B1(_00279_),
    .X(_00280_));
 sky130_fd_sc_hd__nand3_1 _06506_ (.A(net116),
    .B(net59),
    .C(net58),
    .Y(_00281_));
 sky130_fd_sc_hd__a311oi_4 _06507_ (.A1(net118),
    .A2(_00847_),
    .A3(_00000_),
    .B1(_00155_),
    .C1(_00330_),
    .Y(_00282_));
 sky130_fd_sc_hd__a311o_2 _06508_ (.A1(net118),
    .A2(_00847_),
    .A3(_00000_),
    .B1(_00155_),
    .C1(_00330_),
    .X(_00283_));
 sky130_fd_sc_hd__nand2_2 _06509_ (.A(net14),
    .B(net60),
    .Y(_00284_));
 sky130_fd_sc_hd__a22oi_4 _06510_ (.A1(net15),
    .A2(net59),
    .B1(net116),
    .B2(net58),
    .Y(_00285_));
 sky130_fd_sc_hd__nand4b_4 _06511_ (.A_N(_00285_),
    .B(net14),
    .C(_00283_),
    .D(net60),
    .Y(_00287_));
 sky130_fd_sc_hd__o22ai_2 _06512_ (.A1(_00264_),
    .A2(_00281_),
    .B1(_00284_),
    .B2(_00285_),
    .Y(_00288_));
 sky130_fd_sc_hd__o2bb2a_1 _06513_ (.A1_N(_00148_),
    .A2_N(_00149_),
    .B1(_00220_),
    .B2(_00396_),
    .X(_00289_));
 sky130_fd_sc_hd__a22o_1 _06514_ (.A1(net11),
    .A2(net63),
    .B1(_00148_),
    .B2(_00149_),
    .X(_00290_));
 sky130_fd_sc_hd__nor2_1 _06515_ (.A(_00150_),
    .B(_00289_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _06516_ (.A(_00151_),
    .B(_00290_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_2 _06517_ (.A(_00288_),
    .B(_00291_),
    .Y(_00293_));
 sky130_fd_sc_hd__o311a_1 _06518_ (.A1(_00242_),
    .A2(_00352_),
    .A3(_00285_),
    .B1(_00292_),
    .C1(_00283_),
    .X(_00294_));
 sky130_fd_sc_hd__o211ai_2 _06519_ (.A1(_00284_),
    .A2(_00285_),
    .B1(_00292_),
    .C1(_00283_),
    .Y(_00295_));
 sky130_fd_sc_hd__o21ai_1 _06520_ (.A1(_00150_),
    .A2(_00289_),
    .B1(_00288_),
    .Y(_00296_));
 sky130_fd_sc_hd__o211ai_2 _06521_ (.A1(_00284_),
    .A2(_00285_),
    .B1(_00283_),
    .C1(_00291_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand3b_2 _06522_ (.A_N(_00280_),
    .B(_00293_),
    .C(_00295_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand3_2 _06523_ (.A(_00296_),
    .B(_00298_),
    .C(_00280_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand4_1 _06524_ (.A(_00274_),
    .B(_00279_),
    .C(_00293_),
    .D(_00295_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand3b_1 _06525_ (.A_N(_00280_),
    .B(_00296_),
    .C(_00298_),
    .Y(_00302_));
 sky130_fd_sc_hd__o22a_1 _06526_ (.A1(_00264_),
    .A2(_00352_),
    .B1(_00363_),
    .B2(_00869_),
    .X(_00303_));
 sky130_fd_sc_hd__a21oi_2 _06527_ (.A1(_00144_),
    .A2(_00153_),
    .B1(_00303_),
    .Y(_00304_));
 sky130_fd_sc_hd__a31o_1 _06528_ (.A1(net15),
    .A2(net59),
    .A3(_00144_),
    .B1(_00303_),
    .X(_00305_));
 sky130_fd_sc_hd__and3_1 _06529_ (.A(_00299_),
    .B(_00300_),
    .C(_00304_),
    .X(_00306_));
 sky130_fd_sc_hd__nand3_2 _06530_ (.A(_00299_),
    .B(_00300_),
    .C(_00304_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand3_4 _06531_ (.A(_00306_),
    .B(_00272_),
    .C(_00167_),
    .Y(_00309_));
 sky130_fd_sc_hd__a32o_1 _06532_ (.A1(_00299_),
    .A2(_00300_),
    .A3(_00304_),
    .B1(_00272_),
    .B2(_00167_),
    .X(_00310_));
 sky130_fd_sc_hd__nand2_2 _06533_ (.A(net8),
    .B(net34),
    .Y(_00311_));
 sky130_fd_sc_hd__nand4_1 _06534_ (.A(net9),
    .B(net8),
    .C(net64),
    .D(net34),
    .Y(_00312_));
 sky130_fd_sc_hd__a22o_1 _06535_ (.A1(net9),
    .A2(net64),
    .B1(net34),
    .B2(net8),
    .X(_00313_));
 sky130_fd_sc_hd__nand3_1 _06536_ (.A(_00311_),
    .B(net64),
    .C(net9),
    .Y(_00314_));
 sky130_fd_sc_hd__nand3_1 _06537_ (.A(_00171_),
    .B(net34),
    .C(net8),
    .Y(_00315_));
 sky130_fd_sc_hd__nand4_2 _06538_ (.A(_00313_),
    .B(net35),
    .C(net7),
    .D(_00312_),
    .Y(_00316_));
 sky130_fd_sc_hd__o21ai_1 _06539_ (.A1(_00171_),
    .A2(_00311_),
    .B1(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__o22ai_2 _06540_ (.A1(_00209_),
    .A2(_00407_),
    .B1(_00172_),
    .B2(_00173_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand3_2 _06541_ (.A(_00175_),
    .B(_00317_),
    .C(_00318_),
    .Y(_00320_));
 sky130_fd_sc_hd__a22o_1 _06542_ (.A1(net5),
    .A2(net38),
    .B1(_00203_),
    .B2(_00204_),
    .X(_00321_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(_00205_),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__a21o_1 _06544_ (.A1(_00175_),
    .A2(_00318_),
    .B1(_00317_),
    .X(_00323_));
 sky130_fd_sc_hd__nand4_1 _06545_ (.A(_00205_),
    .B(_00320_),
    .C(_00321_),
    .D(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(_00320_),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__a22oi_2 _06547_ (.A1(_00076_),
    .A2(_00181_),
    .B1(_00183_),
    .B2(_00180_),
    .Y(_00326_));
 sky130_fd_sc_hd__a21oi_1 _06548_ (.A1(_00180_),
    .A2(_00183_),
    .B1(_00182_),
    .Y(_00327_));
 sky130_fd_sc_hd__and3_1 _06549_ (.A(_00180_),
    .B(_00182_),
    .C(_00183_),
    .X(_00328_));
 sky130_fd_sc_hd__o2bb2ai_2 _06550_ (.A1_N(_00293_),
    .A2_N(_00299_),
    .B1(_00327_),
    .B2(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__o221ai_4 _06551_ (.A1(_00280_),
    .A2(_00294_),
    .B1(_00326_),
    .B2(_00184_),
    .C1(_00293_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand3_2 _06552_ (.A(_00325_),
    .B(_00329_),
    .C(_00331_),
    .Y(_00332_));
 sky130_fd_sc_hd__a21o_1 _06553_ (.A1(_00329_),
    .A2(_00331_),
    .B1(_00325_),
    .X(_00333_));
 sky130_fd_sc_hd__nand4_4 _06554_ (.A(_00309_),
    .B(_00310_),
    .C(_00332_),
    .D(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__a22oi_4 _06555_ (.A1(_00169_),
    .A2(_00170_),
    .B1(_00195_),
    .B2(_00196_),
    .Y(_00335_));
 sky130_fd_sc_hd__a211oi_1 _06556_ (.A1(_00309_),
    .A2(_00334_),
    .B1(_00335_),
    .C1(_00197_),
    .Y(_00336_));
 sky130_fd_sc_hd__a211o_1 _06557_ (.A1(_00309_),
    .A2(_00334_),
    .B1(_00335_),
    .C1(_00197_),
    .X(_00337_));
 sky130_fd_sc_hd__o2bb2ai_1 _06558_ (.A1_N(_00222_),
    .A2_N(_00223_),
    .B1(_00237_),
    .B2(_00239_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _06559_ (.A(_00241_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand3_1 _06560_ (.A(_00329_),
    .B(_00332_),
    .C(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__a21o_1 _06561_ (.A1(_00329_),
    .A2(_00332_),
    .B1(_00339_),
    .X(_00342_));
 sky130_fd_sc_hd__and4_1 _06562_ (.A(net5),
    .B(net6),
    .C(net37),
    .D(net36),
    .X(_00343_));
 sky130_fd_sc_hd__nand4_1 _06563_ (.A(net5),
    .B(net6),
    .C(net37),
    .D(net36),
    .Y(_00344_));
 sky130_fd_sc_hd__a22o_1 _06564_ (.A1(net5),
    .A2(net37),
    .B1(net36),
    .B2(net6),
    .X(_00345_));
 sky130_fd_sc_hd__and2_1 _06565_ (.A(net4),
    .B(net38),
    .X(_00346_));
 sky130_fd_sc_hd__and3_1 _06566_ (.A(_00344_),
    .B(_00345_),
    .C(_00346_),
    .X(_00347_));
 sky130_fd_sc_hd__a21o_1 _06567_ (.A1(_00345_),
    .A2(_00346_),
    .B1(_00343_),
    .X(_00348_));
 sky130_fd_sc_hd__o211ai_2 _06568_ (.A1(_00143_),
    .A2(_00451_),
    .B1(_00213_),
    .C1(_00214_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand3_1 _06569_ (.A(_00215_),
    .B(_00348_),
    .C(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(net2),
    .B(net40),
    .Y(_00351_));
 sky130_fd_sc_hd__nand4_2 _06571_ (.A(net3),
    .B(net2),
    .C(net39),
    .D(net40),
    .Y(_00353_));
 sky130_fd_sc_hd__a22o_1 _06572_ (.A1(net3),
    .A2(net39),
    .B1(net40),
    .B2(net2),
    .X(_00354_));
 sky130_fd_sc_hd__nand3_1 _06573_ (.A(_00351_),
    .B(net39),
    .C(net3),
    .Y(_00355_));
 sky130_fd_sc_hd__nand3_1 _06574_ (.A(_00210_),
    .B(net40),
    .C(net2),
    .Y(_00356_));
 sky130_fd_sc_hd__nand4_4 _06575_ (.A(_00354_),
    .B(net41),
    .C(net32),
    .D(_00353_),
    .Y(_00357_));
 sky130_fd_sc_hd__o31a_1 _06576_ (.A1(_00132_),
    .A2(_00440_),
    .A3(_00351_),
    .B1(_00357_),
    .X(_00358_));
 sky130_fd_sc_hd__a21oi_1 _06577_ (.A1(_00215_),
    .A2(_00349_),
    .B1(_00348_),
    .Y(_00359_));
 sky130_fd_sc_hd__a21o_1 _06578_ (.A1(_00215_),
    .A2(_00349_),
    .B1(_00348_),
    .X(_00360_));
 sky130_fd_sc_hd__o21a_1 _06579_ (.A1(_00358_),
    .A2(_00359_),
    .B1(_00350_),
    .X(_00361_));
 sky130_fd_sc_hd__a21oi_1 _06580_ (.A1(_00208_),
    .A2(_00218_),
    .B1(_00216_),
    .Y(_00362_));
 sky130_fd_sc_hd__and3_1 _06581_ (.A(_00208_),
    .B(_00218_),
    .C(_00216_),
    .X(_00364_));
 sky130_fd_sc_hd__nand3_1 _06582_ (.A(_00208_),
    .B(_00218_),
    .C(_00216_),
    .Y(_00365_));
 sky130_fd_sc_hd__o21bai_1 _06583_ (.A1(_00362_),
    .A2(_00364_),
    .B1_N(_00361_),
    .Y(_00366_));
 sky130_fd_sc_hd__a22o_1 _06584_ (.A1(net30),
    .A2(net46),
    .B1(net47),
    .B2(net29),
    .X(_00367_));
 sky130_fd_sc_hd__nand4_2 _06585_ (.A(net30),
    .B(net29),
    .C(net46),
    .D(net47),
    .Y(_00368_));
 sky130_fd_sc_hd__a22o_1 _06586_ (.A1(_00367_),
    .A2(_00368_),
    .B1(net117),
    .B2(net28),
    .X(_00369_));
 sky130_fd_sc_hd__nand4_2 _06587_ (.A(net117),
    .B(_00367_),
    .C(_00368_),
    .D(net28),
    .Y(_00370_));
 sky130_fd_sc_hd__nand4_2 _06588_ (.A(net32),
    .B(net31),
    .C(net43),
    .D(net42),
    .Y(_00371_));
 sky130_fd_sc_hd__a22o_1 _06589_ (.A1(net31),
    .A2(net43),
    .B1(net42),
    .B2(net32),
    .X(_00372_));
 sky130_fd_sc_hd__nand4_2 _06590_ (.A(_00372_),
    .B(net45),
    .C(net30),
    .D(_00371_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _06591_ (.A(_00371_),
    .B(_00373_),
    .Y(_00375_));
 sky130_fd_sc_hd__a22o_1 _06592_ (.A1(net31),
    .A2(net45),
    .B1(_00229_),
    .B2(_00230_),
    .X(_00376_));
 sky130_fd_sc_hd__a21o_1 _06593_ (.A1(_00232_),
    .A2(_00376_),
    .B1(_00375_),
    .X(_00377_));
 sky130_fd_sc_hd__nand3_2 _06594_ (.A(_00232_),
    .B(_00375_),
    .C(_00376_),
    .Y(_00378_));
 sky130_fd_sc_hd__a22o_1 _06595_ (.A1(_00369_),
    .A2(_00370_),
    .B1(_00377_),
    .B2(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__nand4_2 _06596_ (.A(_00369_),
    .B(_00370_),
    .C(_00377_),
    .D(_00378_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand3b_1 _06597_ (.A_N(_00362_),
    .B(_00365_),
    .C(_00361_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand4_1 _06598_ (.A(_00366_),
    .B(_00379_),
    .C(_00380_),
    .D(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__nand2_1 _06599_ (.A(_00366_),
    .B(_00382_),
    .Y(_00383_));
 sky130_fd_sc_hd__nand3_1 _06600_ (.A(_00340_),
    .B(_00342_),
    .C(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__a21o_1 _06601_ (.A1(_00340_),
    .A2(_00342_),
    .B1(_00383_),
    .X(_00386_));
 sky130_fd_sc_hd__o211ai_2 _06602_ (.A1(_00197_),
    .A2(_00335_),
    .B1(_00334_),
    .C1(_00309_),
    .Y(_00387_));
 sky130_fd_sc_hd__and4_1 _06603_ (.A(_00337_),
    .B(_00384_),
    .C(_00386_),
    .D(_00387_),
    .X(_00388_));
 sky130_fd_sc_hd__a31o_1 _06604_ (.A1(_00384_),
    .A2(_00386_),
    .A3(_00387_),
    .B1(_00336_),
    .X(_00389_));
 sky130_fd_sc_hd__xor2_1 _06605_ (.A(_00202_),
    .B(_00249_),
    .X(_00390_));
 sky130_fd_sc_hd__o21a_1 _06606_ (.A1(_00336_),
    .A2(_00388_),
    .B1(_00390_),
    .X(_00391_));
 sky130_fd_sc_hd__nand2_1 _06607_ (.A(_00225_),
    .B(_00227_),
    .Y(_00392_));
 sky130_fd_sc_hd__o21a_1 _06608_ (.A1(_00228_),
    .A2(_00236_),
    .B1(_00235_),
    .X(_00393_));
 sky130_fd_sc_hd__and2_1 _06609_ (.A(_00342_),
    .B(_00384_),
    .X(_00394_));
 sky130_fd_sc_hd__xnor2_1 _06610_ (.A(_00393_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__a21o_1 _06611_ (.A1(_00225_),
    .A2(_00227_),
    .B1(_00395_),
    .X(_00397_));
 sky130_fd_sc_hd__xnor2_1 _06612_ (.A(_00392_),
    .B(_00395_),
    .Y(_00398_));
 sky130_fd_sc_hd__nor2_1 _06613_ (.A(_00389_),
    .B(_00390_),
    .Y(_00399_));
 sky130_fd_sc_hd__nor2_1 _06614_ (.A(_00391_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__and2_1 _06615_ (.A(_00398_),
    .B(_00400_),
    .X(_00401_));
 sky130_fd_sc_hd__xnor2_1 _06616_ (.A(_00260_),
    .B(_00261_),
    .Y(_00402_));
 sky130_fd_sc_hd__o21a_1 _06617_ (.A1(_00391_),
    .A2(_00401_),
    .B1(_00402_),
    .X(_00403_));
 sky130_fd_sc_hd__o21ai_1 _06618_ (.A1(_00393_),
    .A2(_00394_),
    .B1(_00397_),
    .Y(_00404_));
 sky130_fd_sc_hd__a211oi_1 _06619_ (.A1(_00389_),
    .A2(_00390_),
    .B1(_00401_),
    .C1(_00402_),
    .Y(_00405_));
 sky130_fd_sc_hd__nor2_1 _06620_ (.A(_00403_),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__a21o_1 _06621_ (.A1(_00406_),
    .A2(_00404_),
    .B1(_00403_),
    .X(_00408_));
 sky130_fd_sc_hd__xnor2_1 _06622_ (.A(_00267_),
    .B(_00268_),
    .Y(_00409_));
 sky130_fd_sc_hd__and2b_1 _06623_ (.A_N(_00409_),
    .B(_00408_),
    .X(_00410_));
 sky130_fd_sc_hd__xor2_2 _06624_ (.A(_00408_),
    .B(_00409_),
    .X(_00411_));
 sky130_fd_sc_hd__xor2_1 _06625_ (.A(_00404_),
    .B(_00406_),
    .X(_00412_));
 sky130_fd_sc_hd__inv_2 _06626_ (.A(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_4 _06627_ (.A(net15),
    .B(net44),
    .Y(_00414_));
 sky130_fd_sc_hd__a21oi_2 _06628_ (.A1(net118),
    .A2(_00858_),
    .B1(_00308_),
    .Y(_00415_));
 sky130_fd_sc_hd__a21oi_1 _06629_ (.A1(net118),
    .A2(_00858_),
    .B1(_00414_),
    .Y(_00416_));
 sky130_fd_sc_hd__and4_2 _06630_ (.A(net116),
    .B(net55),
    .C(net44),
    .D(net15),
    .X(_00417_));
 sky130_fd_sc_hd__o211ai_2 _06631_ (.A1(_00264_),
    .A2(_00308_),
    .B1(net55),
    .C1(net116),
    .Y(_00419_));
 sky130_fd_sc_hd__and2_1 _06632_ (.A(net13),
    .B(net60),
    .X(_00420_));
 sky130_fd_sc_hd__nand2_1 _06633_ (.A(net14),
    .B(net58),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _06634_ (.A(net15),
    .B(net58),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _06635_ (.A(net14),
    .B(net59),
    .Y(_00423_));
 sky130_fd_sc_hd__a22o_1 _06636_ (.A1(net15),
    .A2(net58),
    .B1(net59),
    .B2(net14),
    .X(_00424_));
 sky130_fd_sc_hd__nand3_1 _06637_ (.A(_00423_),
    .B(net58),
    .C(net15),
    .Y(_00425_));
 sky130_fd_sc_hd__nand3_1 _06638_ (.A(_00422_),
    .B(net59),
    .C(net14),
    .Y(_00426_));
 sky130_fd_sc_hd__o2111ai_4 _06639_ (.A1(_00155_),
    .A2(_00421_),
    .B1(net13),
    .C1(net60),
    .D1(_00424_),
    .Y(_00427_));
 sky130_fd_sc_hd__o211ai_4 _06640_ (.A1(_00253_),
    .A2(_00352_),
    .B1(_00425_),
    .C1(_00426_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_2 _06641_ (.A(_00427_),
    .B(_00428_),
    .Y(_00430_));
 sky130_fd_sc_hd__nor2_4 _06642_ (.A(_00419_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__a211oi_2 _06643_ (.A1(_00414_),
    .A2(_00430_),
    .B1(_00341_),
    .C1(_00869_),
    .Y(_00432_));
 sky130_fd_sc_hd__o22a_2 _06644_ (.A1(_00242_),
    .A2(_00352_),
    .B1(_00282_),
    .B2(_00285_),
    .X(_00433_));
 sky130_fd_sc_hd__o21ai_2 _06645_ (.A1(_00282_),
    .A2(_00285_),
    .B1(_00284_),
    .Y(_00434_));
 sky130_fd_sc_hd__o21ai_4 _06646_ (.A1(_00417_),
    .A2(_00431_),
    .B1(_00287_),
    .Y(_00435_));
 sky130_fd_sc_hd__o211ai_4 _06647_ (.A1(_00417_),
    .A2(_00431_),
    .B1(_00434_),
    .C1(_00287_),
    .Y(_00436_));
 sky130_fd_sc_hd__a21oi_2 _06648_ (.A1(_00287_),
    .A2(_00434_),
    .B1(_00432_),
    .Y(_00437_));
 sky130_fd_sc_hd__a21o_2 _06649_ (.A1(_00287_),
    .A2(_00434_),
    .B1(_00432_),
    .X(_00438_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(net10),
    .B(net62),
    .Y(_00439_));
 sky130_fd_sc_hd__nand4_1 _06651_ (.A(net11),
    .B(net10),
    .C(net62),
    .D(net61),
    .Y(_00441_));
 sky130_fd_sc_hd__a22o_1 _06652_ (.A1(net10),
    .A2(net62),
    .B1(net61),
    .B2(net11),
    .X(_00442_));
 sky130_fd_sc_hd__nand4_2 _06653_ (.A(_00442_),
    .B(net63),
    .C(net9),
    .D(_00441_),
    .Y(_00443_));
 sky130_fd_sc_hd__o31a_1 _06654_ (.A1(_00220_),
    .A2(_00385_),
    .A3(_00439_),
    .B1(_00443_),
    .X(_00444_));
 sky130_fd_sc_hd__o2bb2ai_2 _06655_ (.A1_N(_00420_),
    .A2_N(_00424_),
    .B1(_00421_),
    .B2(_00155_),
    .Y(_00445_));
 sky130_fd_sc_hd__o211ai_2 _06656_ (.A1(_00231_),
    .A2(_00396_),
    .B1(_00277_),
    .C1(_00278_),
    .Y(_00446_));
 sky130_fd_sc_hd__a21oi_1 _06657_ (.A1(_00279_),
    .A2(_00446_),
    .B1(_00445_),
    .Y(_00447_));
 sky130_fd_sc_hd__a21o_1 _06658_ (.A1(_00279_),
    .A2(_00446_),
    .B1(_00445_),
    .X(_00448_));
 sky130_fd_sc_hd__nand3_2 _06659_ (.A(_00279_),
    .B(_00445_),
    .C(_00446_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand3b_2 _06660_ (.A_N(_00444_),
    .B(_00448_),
    .C(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__a21bo_1 _06661_ (.A1(_00448_),
    .A2(_00449_),
    .B1_N(_00444_),
    .X(_00452_));
 sky130_fd_sc_hd__nand2_2 _06662_ (.A(_00450_),
    .B(_00452_),
    .Y(_00453_));
 sky130_fd_sc_hd__o2111ai_4 _06663_ (.A1(_00435_),
    .A2(_00433_),
    .B1(_00450_),
    .C1(_00438_),
    .D1(_00452_),
    .Y(_00454_));
 sky130_fd_sc_hd__o22ai_2 _06664_ (.A1(_00433_),
    .A2(_00435_),
    .B1(_00437_),
    .B2(_00453_),
    .Y(_00455_));
 sky130_fd_sc_hd__a21oi_1 _06665_ (.A1(_00299_),
    .A2(_00300_),
    .B1(_00304_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand3_2 _06666_ (.A(_00301_),
    .B(_00302_),
    .C(_00305_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand3_2 _06667_ (.A(_00307_),
    .B(_00455_),
    .C(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__a21o_1 _06668_ (.A1(_00307_),
    .A2(_00457_),
    .B1(_00455_),
    .X(_00459_));
 sky130_fd_sc_hd__o2bb2ai_1 _06669_ (.A1_N(_00436_),
    .A2_N(_00454_),
    .B1(_00456_),
    .B2(_00306_),
    .Y(_00460_));
 sky130_fd_sc_hd__o2111ai_2 _06670_ (.A1(_00453_),
    .A2(_00437_),
    .B1(_00436_),
    .C1(_00307_),
    .D1(_00457_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_2 _06671_ (.A(net7),
    .B(net64),
    .Y(_00463_));
 sky130_fd_sc_hd__and4_1 _06672_ (.A(net7),
    .B(net8),
    .C(net64),
    .D(net34),
    .X(_00464_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(net6),
    .B(net35),
    .Y(_00465_));
 sky130_fd_sc_hd__a22oi_4 _06674_ (.A1(net8),
    .A2(net64),
    .B1(net34),
    .B2(net7),
    .Y(_00466_));
 sky130_fd_sc_hd__a22o_1 _06675_ (.A1(net8),
    .A2(net64),
    .B1(net34),
    .B2(net7),
    .X(_00467_));
 sky130_fd_sc_hd__o2111ai_4 _06676_ (.A1(_00311_),
    .A2(_00463_),
    .B1(net6),
    .C1(net35),
    .D1(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__o22ai_4 _06677_ (.A1(_00311_),
    .A2(_00463_),
    .B1(_00465_),
    .B2(_00466_),
    .Y(_00469_));
 sky130_fd_sc_hd__o211ai_2 _06678_ (.A1(_00176_),
    .A2(_00407_),
    .B1(_00314_),
    .C1(_00315_),
    .Y(_00470_));
 sky130_fd_sc_hd__and3_1 _06679_ (.A(_00316_),
    .B(_00469_),
    .C(_00470_),
    .X(_00471_));
 sky130_fd_sc_hd__nand3_1 _06680_ (.A(_00316_),
    .B(_00469_),
    .C(_00470_),
    .Y(_00472_));
 sky130_fd_sc_hd__a22oi_2 _06681_ (.A1(net4),
    .A2(net38),
    .B1(_00344_),
    .B2(_00345_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _06682_ (.A(_00347_),
    .B(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__a21oi_1 _06683_ (.A1(_00316_),
    .A2(_00470_),
    .B1(_00469_),
    .Y(_00476_));
 sky130_fd_sc_hd__a21o_1 _06684_ (.A1(_00316_),
    .A2(_00470_),
    .B1(_00469_),
    .X(_00477_));
 sky130_fd_sc_hd__and3_1 _06685_ (.A(_00475_),
    .B(_00477_),
    .C(_00472_),
    .X(_00478_));
 sky130_fd_sc_hd__a31o_1 _06686_ (.A1(_00316_),
    .A2(_00469_),
    .A3(_00470_),
    .B1(_00478_),
    .X(_00479_));
 sky130_fd_sc_hd__o21a_1 _06687_ (.A1(_00444_),
    .A2(_00447_),
    .B1(_00449_),
    .X(_00480_));
 sky130_fd_sc_hd__o21ai_1 _06688_ (.A1(_00444_),
    .A2(_00447_),
    .B1(_00449_),
    .Y(_00481_));
 sky130_fd_sc_hd__a22o_1 _06689_ (.A1(_00205_),
    .A2(_00321_),
    .B1(_00323_),
    .B2(_00320_),
    .X(_00482_));
 sky130_fd_sc_hd__a21o_1 _06690_ (.A1(_00320_),
    .A2(_00323_),
    .B1(_00322_),
    .X(_00483_));
 sky130_fd_sc_hd__nand3_1 _06691_ (.A(_00320_),
    .B(_00322_),
    .C(_00323_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand3_2 _06692_ (.A(_00324_),
    .B(_00481_),
    .C(_00482_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand3_2 _06693_ (.A(_00483_),
    .B(_00485_),
    .C(_00480_),
    .Y(_00487_));
 sky130_fd_sc_hd__o211a_1 _06694_ (.A1(_00471_),
    .A2(_00478_),
    .B1(_00486_),
    .C1(_00487_),
    .X(_00488_));
 sky130_fd_sc_hd__o211ai_2 _06695_ (.A1(_00471_),
    .A2(_00478_),
    .B1(_00486_),
    .C1(_00487_),
    .Y(_00489_));
 sky130_fd_sc_hd__a21oi_1 _06696_ (.A1(_00486_),
    .A2(_00487_),
    .B1(_00479_),
    .Y(_00490_));
 sky130_fd_sc_hd__a211o_1 _06697_ (.A1(_00486_),
    .A2(_00487_),
    .B1(_00471_),
    .C1(_00478_),
    .X(_00491_));
 sky130_fd_sc_hd__nand4_4 _06698_ (.A(_00458_),
    .B(_00459_),
    .C(_00489_),
    .D(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(_00458_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__a22o_1 _06700_ (.A1(_00309_),
    .A2(_00310_),
    .B1(_00332_),
    .B2(_00333_),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _06701_ (.A1(_00458_),
    .A2(_00492_),
    .B1(_00494_),
    .B2(_00334_),
    .X(_00496_));
 sky130_fd_sc_hd__nand4_1 _06702_ (.A(_00334_),
    .B(_00458_),
    .C(_00492_),
    .D(_00494_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand4_2 _06703_ (.A(net5),
    .B(net4),
    .C(net37),
    .D(net36),
    .Y(_00498_));
 sky130_fd_sc_hd__a22oi_1 _06704_ (.A1(net4),
    .A2(net37),
    .B1(net36),
    .B2(net5),
    .Y(_00499_));
 sky130_fd_sc_hd__a22o_1 _06705_ (.A1(net4),
    .A2(net37),
    .B1(net36),
    .B2(net5),
    .X(_00500_));
 sky130_fd_sc_hd__nand2_1 _06706_ (.A(net3),
    .B(net38),
    .Y(_00501_));
 sky130_fd_sc_hd__nand4_4 _06707_ (.A(_00500_),
    .B(net38),
    .C(net3),
    .D(_00498_),
    .Y(_00502_));
 sky130_fd_sc_hd__o21ai_1 _06708_ (.A1(_00501_),
    .A2(_00499_),
    .B1(_00498_),
    .Y(_00503_));
 sky130_fd_sc_hd__o211ai_2 _06709_ (.A1(_00110_),
    .A2(_00451_),
    .B1(_00355_),
    .C1(_00356_),
    .Y(_00504_));
 sky130_fd_sc_hd__and3_1 _06710_ (.A(_00357_),
    .B(_00503_),
    .C(_00504_),
    .X(_00505_));
 sky130_fd_sc_hd__nand3_1 _06711_ (.A(_00357_),
    .B(_00503_),
    .C(_00504_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand4_4 _06712_ (.A(net32),
    .B(net2),
    .C(net39),
    .D(net40),
    .Y(_00508_));
 sky130_fd_sc_hd__a22o_1 _06713_ (.A1(net2),
    .A2(net39),
    .B1(net40),
    .B2(net32),
    .X(_00509_));
 sky130_fd_sc_hd__nand3_2 _06714_ (.A(_00509_),
    .B(net41),
    .C(_00508_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand4_2 _06715_ (.A(_00509_),
    .B(net41),
    .C(net31),
    .D(_00508_),
    .Y(_00511_));
 sky130_fd_sc_hd__o31a_1 _06716_ (.A1(_00110_),
    .A2(_00440_),
    .A3(_00351_),
    .B1(_00511_),
    .X(_00512_));
 sky130_fd_sc_hd__a21oi_1 _06717_ (.A1(_00357_),
    .A2(_00504_),
    .B1(_00503_),
    .Y(_00513_));
 sky130_fd_sc_hd__a21o_1 _06718_ (.A1(_00357_),
    .A2(_00504_),
    .B1(_00503_),
    .X(_00514_));
 sky130_fd_sc_hd__a211oi_1 _06719_ (.A1(_00508_),
    .A2(_00511_),
    .B1(_00513_),
    .C1(_00505_),
    .Y(_00515_));
 sky130_fd_sc_hd__o21a_1 _06720_ (.A1(_00512_),
    .A2(_00513_),
    .B1(_00507_),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _06721_ (.A1(_00353_),
    .A2(_00357_),
    .B1(_00360_),
    .B2(_00350_),
    .X(_00518_));
 sky130_fd_sc_hd__nand3_1 _06722_ (.A(_00350_),
    .B(_00360_),
    .C(_00358_),
    .Y(_00519_));
 sky130_fd_sc_hd__a21o_1 _06723_ (.A1(_00518_),
    .A2(_00519_),
    .B1(_00516_),
    .X(_00520_));
 sky130_fd_sc_hd__a22o_1 _06724_ (.A1(net29),
    .A2(net46),
    .B1(net47),
    .B2(net28),
    .X(_00521_));
 sky130_fd_sc_hd__nand4_2 _06725_ (.A(net28),
    .B(net29),
    .C(net46),
    .D(net47),
    .Y(_00522_));
 sky130_fd_sc_hd__a22o_1 _06726_ (.A1(_00521_),
    .A2(_00522_),
    .B1(net117),
    .B2(net27),
    .X(_00523_));
 sky130_fd_sc_hd__nand4_2 _06727_ (.A(net117),
    .B(_00521_),
    .C(_00522_),
    .D(net27),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_2 _06728_ (.A(net30),
    .B(net43),
    .Y(_00525_));
 sky130_fd_sc_hd__and4_1 _06729_ (.A(net30),
    .B(net31),
    .C(net43),
    .D(net42),
    .X(_00526_));
 sky130_fd_sc_hd__nand4_2 _06730_ (.A(net30),
    .B(net31),
    .C(net43),
    .D(net42),
    .Y(_00527_));
 sky130_fd_sc_hd__a22o_1 _06731_ (.A1(net30),
    .A2(net43),
    .B1(net42),
    .B2(net31),
    .X(_00529_));
 sky130_fd_sc_hd__and4_2 _06732_ (.A(_00529_),
    .B(net45),
    .C(net29),
    .D(_00527_),
    .X(_00530_));
 sky130_fd_sc_hd__a22o_1 _06733_ (.A1(net30),
    .A2(net45),
    .B1(_00371_),
    .B2(_00372_),
    .X(_00531_));
 sky130_fd_sc_hd__a211o_1 _06734_ (.A1(_00373_),
    .A2(_00531_),
    .B1(_00530_),
    .C1(_00526_),
    .X(_00532_));
 sky130_fd_sc_hd__o211ai_4 _06735_ (.A1(_00526_),
    .A2(_00530_),
    .B1(_00531_),
    .C1(_00373_),
    .Y(_00533_));
 sky130_fd_sc_hd__a22o_1 _06736_ (.A1(_00523_),
    .A2(_00524_),
    .B1(_00532_),
    .B2(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__nand4_2 _06737_ (.A(_00523_),
    .B(_00524_),
    .C(_00532_),
    .D(_00533_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand3_1 _06738_ (.A(_00516_),
    .B(_00518_),
    .C(_00519_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand4_2 _06739_ (.A(_00520_),
    .B(_00534_),
    .C(_00535_),
    .D(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(_00520_),
    .B(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _06741_ (.A(_00486_),
    .B(_00489_),
    .Y(_00540_));
 sky130_fd_sc_hd__a22o_1 _06742_ (.A1(_00379_),
    .A2(_00380_),
    .B1(_00381_),
    .B2(_00366_),
    .X(_00541_));
 sky130_fd_sc_hd__nand3_1 _06743_ (.A(_00382_),
    .B(_00540_),
    .C(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__a21o_1 _06744_ (.A1(_00382_),
    .A2(_00541_),
    .B1(_00540_),
    .X(_00543_));
 sky130_fd_sc_hd__a22o_1 _06745_ (.A1(_00520_),
    .A2(_00537_),
    .B1(_00542_),
    .B2(_00543_),
    .X(_00544_));
 sky130_fd_sc_hd__nand4_1 _06746_ (.A(_00520_),
    .B(_00537_),
    .C(_00542_),
    .D(_00543_),
    .Y(_00545_));
 sky130_fd_sc_hd__a22oi_2 _06747_ (.A1(_00496_),
    .A2(_00497_),
    .B1(_00544_),
    .B2(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__a31o_1 _06748_ (.A1(_00334_),
    .A2(_00493_),
    .A3(_00494_),
    .B1(_00546_),
    .X(_00547_));
 sky130_fd_sc_hd__a22oi_1 _06749_ (.A1(_00384_),
    .A2(_00386_),
    .B1(_00387_),
    .B2(_00337_),
    .Y(_00548_));
 sky130_fd_sc_hd__nor2_1 _06750_ (.A(_00388_),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(_00549_),
    .B(_00547_),
    .Y(_00551_));
 sky130_fd_sc_hd__xnor2_1 _06752_ (.A(_00547_),
    .B(_00549_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_2 _06753_ (.A(_00368_),
    .B(_00370_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_2 _06754_ (.A(_00378_),
    .B(_00380_),
    .Y(_00554_));
 sky130_fd_sc_hd__a21bo_2 _06755_ (.A1(_00538_),
    .A2(_00543_),
    .B1_N(_00542_),
    .X(_00555_));
 sky130_fd_sc_hd__xor2_2 _06756_ (.A(_00554_),
    .B(_00555_),
    .X(_00556_));
 sky130_fd_sc_hd__xnor2_1 _06757_ (.A(_00553_),
    .B(_00556_),
    .Y(_00557_));
 sky130_fd_sc_hd__or2_1 _06758_ (.A(_00552_),
    .B(_00557_),
    .X(_00558_));
 sky130_fd_sc_hd__nor2_1 _06759_ (.A(_00398_),
    .B(_00400_),
    .Y(_00559_));
 sky130_fd_sc_hd__o221a_1 _06760_ (.A1(_00552_),
    .A2(_00557_),
    .B1(_00559_),
    .B2(_00401_),
    .C1(_00551_),
    .X(_00560_));
 sky130_fd_sc_hd__a211o_1 _06761_ (.A1(_00551_),
    .A2(_00558_),
    .B1(_00559_),
    .C1(_00401_),
    .X(_00562_));
 sky130_fd_sc_hd__a22oi_1 _06762_ (.A1(_00554_),
    .A2(_00555_),
    .B1(_00556_),
    .B2(_00553_),
    .Y(_00563_));
 sky130_fd_sc_hd__o21a_1 _06763_ (.A1(_00560_),
    .A2(_00563_),
    .B1(_00562_),
    .X(_00564_));
 sky130_fd_sc_hd__nor2_1 _06764_ (.A(_00413_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _06765_ (.A(_00552_),
    .B(_00557_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _06766_ (.A(_00558_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__a32oi_4 _06767_ (.A1(net116),
    .A2(_00414_),
    .A3(net55),
    .B1(_00427_),
    .B2(_00428_),
    .Y(_00568_));
 sky130_fd_sc_hd__and4_1 _06768_ (.A(net116),
    .B(_00414_),
    .C(_00430_),
    .D(net55),
    .X(_00569_));
 sky130_fd_sc_hd__and3_1 _06769_ (.A(_00419_),
    .B(_00427_),
    .C(_00428_),
    .X(_00570_));
 sky130_fd_sc_hd__a22oi_4 _06770_ (.A1(net15),
    .A2(net55),
    .B1(net116),
    .B2(net44),
    .Y(_00571_));
 sky130_fd_sc_hd__a21oi_1 _06771_ (.A1(net55),
    .A2(_00416_),
    .B1(_00571_),
    .Y(_00573_));
 sky130_fd_sc_hd__a21o_1 _06772_ (.A1(net55),
    .A2(_00416_),
    .B1(_00571_),
    .X(_00574_));
 sky130_fd_sc_hd__nor2_2 _06773_ (.A(_00264_),
    .B(_00319_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(net15),
    .B(net33),
    .Y(_00576_));
 sky130_fd_sc_hd__nand4_2 _06775_ (.A(net116),
    .B(net33),
    .C(net44),
    .D(net15),
    .Y(_00577_));
 sky130_fd_sc_hd__nor2_1 _06776_ (.A(_00242_),
    .B(_00341_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(net14),
    .B(net55),
    .Y(_00579_));
 sky130_fd_sc_hd__a22oi_4 _06778_ (.A1(net15),
    .A2(net44),
    .B1(net116),
    .B2(net33),
    .Y(_00580_));
 sky130_fd_sc_hd__o2bb2ai_4 _06779_ (.A1_N(net33),
    .A2_N(net116),
    .B1(_00264_),
    .B2(_00308_),
    .Y(_00581_));
 sky130_fd_sc_hd__a211oi_4 _06780_ (.A1(_00415_),
    .A2(_00575_),
    .B1(_00579_),
    .C1(_00580_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand4_2 _06781_ (.A(_00581_),
    .B(net55),
    .C(net14),
    .D(_00577_),
    .Y(_00584_));
 sky130_fd_sc_hd__a22oi_4 _06782_ (.A1(_00415_),
    .A2(_00575_),
    .B1(_00581_),
    .B2(_00578_),
    .Y(_00585_));
 sky130_fd_sc_hd__o21ai_1 _06783_ (.A1(_00579_),
    .A2(_00580_),
    .B1(_00577_),
    .Y(_00586_));
 sky130_fd_sc_hd__o21ai_4 _06784_ (.A1(_00417_),
    .A2(_00571_),
    .B1(_00585_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_2 _06785_ (.A(_00586_),
    .B(_00573_),
    .Y(_00588_));
 sky130_fd_sc_hd__and4_2 _06786_ (.A(net14),
    .B(net13),
    .C(net58),
    .D(net59),
    .X(_00589_));
 sky130_fd_sc_hd__o22a_1 _06787_ (.A1(_00242_),
    .A2(_00330_),
    .B1(_00363_),
    .B2(_00253_),
    .X(_00590_));
 sky130_fd_sc_hd__a22o_1 _06788_ (.A1(net14),
    .A2(net58),
    .B1(net59),
    .B2(net13),
    .X(_00591_));
 sky130_fd_sc_hd__and4b_2 _06789_ (.A_N(_00589_),
    .B(_00591_),
    .C(net11),
    .D(net60),
    .X(_00592_));
 sky130_fd_sc_hd__o22a_2 _06790_ (.A1(_00220_),
    .A2(_00352_),
    .B1(_00589_),
    .B2(_00590_),
    .X(_00593_));
 sky130_fd_sc_hd__a211oi_4 _06791_ (.A1(net11),
    .A2(net60),
    .B1(_00589_),
    .C1(_00590_),
    .Y(_00595_));
 sky130_fd_sc_hd__o211a_2 _06792_ (.A1(_00589_),
    .A2(_00590_),
    .B1(net11),
    .C1(net60),
    .X(_00596_));
 sky130_fd_sc_hd__o22ai_2 _06793_ (.A1(_00592_),
    .A2(_00593_),
    .B1(_00574_),
    .B2(_00585_),
    .Y(_00597_));
 sky130_fd_sc_hd__o22ai_2 _06794_ (.A1(_00595_),
    .A2(_00596_),
    .B1(_00573_),
    .B2(_00586_),
    .Y(_00598_));
 sky130_fd_sc_hd__o211ai_4 _06795_ (.A1(_00569_),
    .A2(_00570_),
    .B1(_00587_),
    .C1(_00597_),
    .Y(_00599_));
 sky130_fd_sc_hd__o211ai_4 _06796_ (.A1(_00431_),
    .A2(_00568_),
    .B1(_00588_),
    .C1(_00598_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_2 _06797_ (.A(net9),
    .B(net61),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _06798_ (.A(net9),
    .B(net62),
    .Y(_00602_));
 sky130_fd_sc_hd__and4_1 _06799_ (.A(net9),
    .B(net10),
    .C(net62),
    .D(net61),
    .X(_00603_));
 sky130_fd_sc_hd__a22oi_1 _06800_ (.A1(net9),
    .A2(net62),
    .B1(net61),
    .B2(net10),
    .Y(_00604_));
 sky130_fd_sc_hd__a22o_1 _06801_ (.A1(net9),
    .A2(net62),
    .B1(net61),
    .B2(net10),
    .X(_00606_));
 sky130_fd_sc_hd__o2111a_1 _06802_ (.A1(_00439_),
    .A2(_00601_),
    .B1(net8),
    .C1(net63),
    .D1(_00606_),
    .X(_00607_));
 sky130_fd_sc_hd__o2111ai_4 _06803_ (.A1(_00439_),
    .A2(_00601_),
    .B1(net8),
    .C1(net63),
    .D1(_00606_),
    .Y(_00608_));
 sky130_fd_sc_hd__a31o_1 _06804_ (.A1(_00606_),
    .A2(net63),
    .A3(net8),
    .B1(_00603_),
    .X(_00609_));
 sky130_fd_sc_hd__a31o_1 _06805_ (.A1(_00591_),
    .A2(net60),
    .A3(net11),
    .B1(_00589_),
    .X(_00610_));
 sky130_fd_sc_hd__o2bb2ai_1 _06806_ (.A1_N(_00441_),
    .A2_N(_00442_),
    .B1(_00198_),
    .B2(_00396_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand3_2 _06807_ (.A(_00443_),
    .B(_00610_),
    .C(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__a21o_1 _06808_ (.A1(_00443_),
    .A2(_00611_),
    .B1(_00610_),
    .X(_00613_));
 sky130_fd_sc_hd__o211a_1 _06809_ (.A1(_00603_),
    .A2(_00607_),
    .B1(_00612_),
    .C1(_00613_),
    .X(_00614_));
 sky130_fd_sc_hd__o211ai_2 _06810_ (.A1(_00603_),
    .A2(_00607_),
    .B1(_00612_),
    .C1(_00613_),
    .Y(_00615_));
 sky130_fd_sc_hd__a21oi_1 _06811_ (.A1(_00612_),
    .A2(_00613_),
    .B1(_00609_),
    .Y(_00617_));
 sky130_fd_sc_hd__nor2_1 _06812_ (.A(_00614_),
    .B(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand3_2 _06813_ (.A(_00599_),
    .B(_00600_),
    .C(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__a21boi_1 _06814_ (.A1(_00600_),
    .A2(_00618_),
    .B1_N(_00599_),
    .Y(_00620_));
 sky130_fd_sc_hd__a22o_1 _06815_ (.A1(_00436_),
    .A2(_00438_),
    .B1(_00450_),
    .B2(_00452_),
    .X(_00621_));
 sky130_fd_sc_hd__o211ai_2 _06816_ (.A1(_00435_),
    .A2(_00433_),
    .B1(_00453_),
    .C1(_00438_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21o_1 _06817_ (.A1(_00436_),
    .A2(_00438_),
    .B1(_00453_),
    .X(_00623_));
 sky130_fd_sc_hd__a21oi_1 _06818_ (.A1(_00622_),
    .A2(_00623_),
    .B1(_00620_),
    .Y(_00624_));
 sky130_fd_sc_hd__a22o_1 _06819_ (.A1(_00599_),
    .A2(_00619_),
    .B1(_00622_),
    .B2(_00623_),
    .X(_00625_));
 sky130_fd_sc_hd__nand4_2 _06820_ (.A(net7),
    .B(net6),
    .C(net64),
    .D(net34),
    .Y(_00626_));
 sky130_fd_sc_hd__a22o_1 _06821_ (.A1(net7),
    .A2(net64),
    .B1(net34),
    .B2(net6),
    .X(_00628_));
 sky130_fd_sc_hd__and2_1 _06822_ (.A(net5),
    .B(net35),
    .X(_00629_));
 sky130_fd_sc_hd__nand3_2 _06823_ (.A(_00628_),
    .B(net35),
    .C(_00626_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand4_1 _06824_ (.A(_00628_),
    .B(net35),
    .C(net5),
    .D(_00626_),
    .Y(_00631_));
 sky130_fd_sc_hd__a21bo_1 _06825_ (.A1(_00628_),
    .A2(_00629_),
    .B1_N(_00626_),
    .X(_00632_));
 sky130_fd_sc_hd__o22ai_4 _06826_ (.A1(_00187_),
    .A2(_00407_),
    .B1(_00464_),
    .B2(_00466_),
    .Y(_00633_));
 sky130_fd_sc_hd__and3_1 _06827_ (.A(_00468_),
    .B(_00632_),
    .C(_00633_),
    .X(_00634_));
 sky130_fd_sc_hd__nand3_4 _06828_ (.A(_00468_),
    .B(_00632_),
    .C(_00633_),
    .Y(_00635_));
 sky130_fd_sc_hd__a22o_2 _06829_ (.A1(net3),
    .A2(net38),
    .B1(_00498_),
    .B2(_00500_),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(_00502_),
    .B(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__a21oi_1 _06831_ (.A1(_00468_),
    .A2(_00633_),
    .B1(_00632_),
    .Y(_00639_));
 sky130_fd_sc_hd__a21o_1 _06832_ (.A1(_00468_),
    .A2(_00633_),
    .B1(_00632_),
    .X(_00640_));
 sky130_fd_sc_hd__nor3_2 _06833_ (.A(_00637_),
    .B(_00639_),
    .C(_00634_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand4_2 _06834_ (.A(_00502_),
    .B(_00635_),
    .C(_00636_),
    .D(_00640_),
    .Y(_00642_));
 sky130_fd_sc_hd__o21a_1 _06835_ (.A1(_00637_),
    .A2(_00639_),
    .B1(_00635_),
    .X(_00643_));
 sky130_fd_sc_hd__o21ai_1 _06836_ (.A1(_00471_),
    .A2(_00476_),
    .B1(_00475_),
    .Y(_00644_));
 sky130_fd_sc_hd__o211ai_1 _06837_ (.A1(_00347_),
    .A2(_00474_),
    .B1(_00477_),
    .C1(_00472_),
    .Y(_00645_));
 sky130_fd_sc_hd__a22o_1 _06838_ (.A1(_00612_),
    .A2(_00615_),
    .B1(_00644_),
    .B2(_00645_),
    .X(_00646_));
 sky130_fd_sc_hd__nand4_1 _06839_ (.A(_00612_),
    .B(_00615_),
    .C(_00644_),
    .D(_00645_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_00646_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__a21o_1 _06841_ (.A1(_00635_),
    .A2(_00642_),
    .B1(_00648_),
    .X(_00650_));
 sky130_fd_sc_hd__a211o_2 _06842_ (.A1(_00646_),
    .A2(_00647_),
    .B1(_00634_),
    .C1(_00641_),
    .X(_00651_));
 sky130_fd_sc_hd__a22o_1 _06843_ (.A1(_00635_),
    .A2(_00642_),
    .B1(_00646_),
    .B2(_00647_),
    .X(_00652_));
 sky130_fd_sc_hd__a311o_1 _06844_ (.A1(_00468_),
    .A2(_00632_),
    .A3(_00633_),
    .B1(_00641_),
    .C1(_00648_),
    .X(_00653_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(_00650_),
    .B(_00651_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand3_2 _06846_ (.A(_00620_),
    .B(_00622_),
    .C(_00623_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand4_1 _06847_ (.A(_00454_),
    .B(_00599_),
    .C(_00619_),
    .D(_00621_),
    .Y(_00656_));
 sky130_fd_sc_hd__a22o_1 _06848_ (.A1(_00599_),
    .A2(_00619_),
    .B1(_00621_),
    .B2(_00454_),
    .X(_00657_));
 sky130_fd_sc_hd__nand4_4 _06849_ (.A(_00625_),
    .B(_00650_),
    .C(_00651_),
    .D(_00655_),
    .Y(_00658_));
 sky130_fd_sc_hd__a31o_1 _06850_ (.A1(_00650_),
    .A2(_00651_),
    .A3(_00655_),
    .B1(_00624_),
    .X(_00659_));
 sky130_fd_sc_hd__o211ai_2 _06851_ (.A1(_00488_),
    .A2(_00490_),
    .B1(_00460_),
    .C1(_00461_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(_00492_),
    .B(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand3_2 _06853_ (.A(_00492_),
    .B(_00659_),
    .C(_00661_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand3_2 _06854_ (.A(_00625_),
    .B(_00658_),
    .C(_00662_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand4_1 _06855_ (.A(net3),
    .B(net4),
    .C(net37),
    .D(net36),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(net3),
    .B(net37),
    .Y(_00666_));
 sky130_fd_sc_hd__a22o_1 _06857_ (.A1(net3),
    .A2(net37),
    .B1(net36),
    .B2(net4),
    .X(_00667_));
 sky130_fd_sc_hd__and2_1 _06858_ (.A(net2),
    .B(net38),
    .X(_00668_));
 sky130_fd_sc_hd__and4_1 _06859_ (.A(_00667_),
    .B(net38),
    .C(net2),
    .D(_00665_),
    .X(_00669_));
 sky130_fd_sc_hd__a21bo_1 _06860_ (.A1(_00667_),
    .A2(_00668_),
    .B1_N(_00665_),
    .X(_00670_));
 sky130_fd_sc_hd__a22o_1 _06861_ (.A1(net31),
    .A2(net41),
    .B1(_00508_),
    .B2(_00509_),
    .X(_00672_));
 sky130_fd_sc_hd__o211a_1 _06862_ (.A1(_00121_),
    .A2(_00510_),
    .B1(_00670_),
    .C1(_00672_),
    .X(_00673_));
 sky130_fd_sc_hd__o211ai_4 _06863_ (.A1(_00121_),
    .A2(_00510_),
    .B1(_00670_),
    .C1(_00672_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(net31),
    .B(net39),
    .Y(_00675_));
 sky130_fd_sc_hd__and4_1 _06865_ (.A(net32),
    .B(net31),
    .C(net39),
    .D(net40),
    .X(_00676_));
 sky130_fd_sc_hd__a22oi_2 _06866_ (.A1(net32),
    .A2(net39),
    .B1(net40),
    .B2(net31),
    .Y(_00677_));
 sky130_fd_sc_hd__a22o_1 _06867_ (.A1(net32),
    .A2(net39),
    .B1(net40),
    .B2(net31),
    .X(_00678_));
 sky130_fd_sc_hd__nand4b_2 _06868_ (.A_N(_00676_),
    .B(_00678_),
    .C(net30),
    .D(net41),
    .Y(_00679_));
 sky130_fd_sc_hd__a31o_1 _06869_ (.A1(_00678_),
    .A2(net41),
    .A3(net30),
    .B1(_00676_),
    .X(_00680_));
 sky130_fd_sc_hd__a21oi_1 _06870_ (.A1(_00511_),
    .A2(_00672_),
    .B1(_00670_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21o_1 _06871_ (.A1(_00511_),
    .A2(_00672_),
    .B1(_00670_),
    .X(_00683_));
 sky130_fd_sc_hd__nand3_2 _06872_ (.A(_00674_),
    .B(_00680_),
    .C(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__a21boi_1 _06873_ (.A1(_00507_),
    .A2(_00514_),
    .B1_N(_00512_),
    .Y(_00685_));
 sky130_fd_sc_hd__a21oi_1 _06874_ (.A1(_00507_),
    .A2(_00514_),
    .B1(_00512_),
    .Y(_00686_));
 sky130_fd_sc_hd__and3_1 _06875_ (.A(_00507_),
    .B(_00514_),
    .C(_00512_),
    .X(_00687_));
 sky130_fd_sc_hd__o2bb2ai_2 _06876_ (.A1_N(_00674_),
    .A2_N(_00684_),
    .B1(_00686_),
    .B2(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__a22o_1 _06877_ (.A1(net28),
    .A2(net46),
    .B1(net47),
    .B2(net27),
    .X(_00689_));
 sky130_fd_sc_hd__nand4_2 _06878_ (.A(net28),
    .B(net27),
    .C(net46),
    .D(net47),
    .Y(_00690_));
 sky130_fd_sc_hd__a22o_1 _06879_ (.A1(_00689_),
    .A2(_00690_),
    .B1(net117),
    .B2(net26),
    .X(_00691_));
 sky130_fd_sc_hd__nand4_2 _06880_ (.A(net117),
    .B(_00689_),
    .C(_00690_),
    .D(net26),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_2 _06881_ (.A(net29),
    .B(net42),
    .Y(_00694_));
 sky130_fd_sc_hd__nand4_1 _06882_ (.A(net30),
    .B(net29),
    .C(net43),
    .D(net42),
    .Y(_00695_));
 sky130_fd_sc_hd__a22o_1 _06883_ (.A1(net29),
    .A2(net43),
    .B1(net42),
    .B2(net30),
    .X(_00696_));
 sky130_fd_sc_hd__o2111ai_4 _06884_ (.A1(_00525_),
    .A2(_00694_),
    .B1(net28),
    .C1(net45),
    .D1(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__a22oi_4 _06885_ (.A1(net29),
    .A2(net45),
    .B1(_00527_),
    .B2(_00529_),
    .Y(_00698_));
 sky130_fd_sc_hd__o221ai_4 _06886_ (.A1(_00525_),
    .A2(_00694_),
    .B1(_00698_),
    .B2(_00530_),
    .C1(_00697_),
    .Y(_00699_));
 sky130_fd_sc_hd__a211o_1 _06887_ (.A1(_00695_),
    .A2(_00697_),
    .B1(_00698_),
    .C1(_00530_),
    .X(_00700_));
 sky130_fd_sc_hd__a22o_1 _06888_ (.A1(_00691_),
    .A2(_00692_),
    .B1(_00699_),
    .B2(_00700_),
    .X(_00701_));
 sky130_fd_sc_hd__nand4_2 _06889_ (.A(_00691_),
    .B(_00692_),
    .C(_00699_),
    .D(_00700_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _06890_ (.A(_00701_),
    .B(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__o211ai_2 _06891_ (.A1(_00515_),
    .A2(_00685_),
    .B1(_00684_),
    .C1(_00674_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand4_1 _06892_ (.A(_00688_),
    .B(_00701_),
    .C(_00702_),
    .D(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _06893_ (.A(_00688_),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__o21ai_2 _06894_ (.A1(_00643_),
    .A2(_00648_),
    .B1(_00646_),
    .Y(_00708_));
 sky130_fd_sc_hd__a22o_1 _06895_ (.A1(_00534_),
    .A2(_00535_),
    .B1(_00536_),
    .B2(_00520_),
    .X(_00709_));
 sky130_fd_sc_hd__nand3_2 _06896_ (.A(_00537_),
    .B(_00708_),
    .C(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__a21o_1 _06897_ (.A1(_00537_),
    .A2(_00709_),
    .B1(_00708_),
    .X(_00711_));
 sky130_fd_sc_hd__nand3_2 _06898_ (.A(_00707_),
    .B(_00710_),
    .C(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__a21o_1 _06899_ (.A1(_00710_),
    .A2(_00711_),
    .B1(_00707_),
    .X(_00713_));
 sky130_fd_sc_hd__nand4_2 _06900_ (.A(_00663_),
    .B(_00664_),
    .C(_00712_),
    .D(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__and4_1 _06901_ (.A(_00496_),
    .B(_00497_),
    .C(_00544_),
    .D(_00545_),
    .X(_00716_));
 sky130_fd_sc_hd__a211oi_1 _06902_ (.A1(_00663_),
    .A2(_00714_),
    .B1(_00716_),
    .C1(_00546_),
    .Y(_00717_));
 sky130_fd_sc_hd__o211a_1 _06903_ (.A1(_00546_),
    .A2(_00716_),
    .B1(_00714_),
    .C1(_00663_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_00522_),
    .B(_00524_),
    .Y(_00719_));
 sky130_fd_sc_hd__a22oi_2 _06905_ (.A1(_00533_),
    .A2(_00535_),
    .B1(_00710_),
    .B2(_00712_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand4_1 _06906_ (.A(_00533_),
    .B(_00535_),
    .C(_00710_),
    .D(_00712_),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _06907_ (.A(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__a211o_1 _06908_ (.A1(_00522_),
    .A2(_00524_),
    .B1(_00720_),
    .C1(_00722_),
    .X(_00723_));
 sky130_fd_sc_hd__o21bai_1 _06909_ (.A1(_00720_),
    .A2(_00722_),
    .B1_N(_00719_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(_00723_),
    .B(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__o21ba_1 _06911_ (.A1(_00718_),
    .A2(_00725_),
    .B1_N(_00717_),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _06912_ (.A(_00727_),
    .B(_00567_),
    .X(_00728_));
 sky130_fd_sc_hd__a21oi_1 _06913_ (.A1(_00719_),
    .A2(_00721_),
    .B1(_00720_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _06914_ (.A(_00567_),
    .B(_00727_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _06915_ (.A(_00728_),
    .B(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__or2_1 _06916_ (.A(_00729_),
    .B(_00731_),
    .X(_00732_));
 sky130_fd_sc_hd__o21a_1 _06917_ (.A1(_00729_),
    .A2(_00731_),
    .B1(_00728_),
    .X(_00733_));
 sky130_fd_sc_hd__and2b_1 _06918_ (.A_N(_00560_),
    .B(_00562_),
    .X(_00734_));
 sky130_fd_sc_hd__a221oi_4 _06919_ (.A1(_00554_),
    .A2(_00555_),
    .B1(_00556_),
    .B2(_00553_),
    .C1(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__and2b_1 _06920_ (.A_N(_00563_),
    .B(_00734_),
    .X(_00736_));
 sky130_fd_sc_hd__or3_1 _06921_ (.A(_00733_),
    .B(_00735_),
    .C(_00736_),
    .X(_00738_));
 sky130_fd_sc_hd__o21ai_1 _06922_ (.A1(_00735_),
    .A2(_00736_),
    .B1(_00733_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_2 _06923_ (.A(_00738_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__nand3_2 _06924_ (.A(_00654_),
    .B(_00656_),
    .C(_00657_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand4_1 _06925_ (.A(_00625_),
    .B(_00652_),
    .C(_00653_),
    .D(_00655_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand4_1 _06926_ (.A(_00650_),
    .B(_00651_),
    .C(_00656_),
    .D(_00657_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_2 _06927_ (.A(net14),
    .B(net33),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_2 _06928_ (.A(net14),
    .B(net44),
    .Y(_00745_));
 sky130_fd_sc_hd__a22o_1 _06929_ (.A1(net14),
    .A2(net44),
    .B1(net33),
    .B2(net15),
    .X(_00746_));
 sky130_fd_sc_hd__nand3_1 _06930_ (.A(_00745_),
    .B(net33),
    .C(net15),
    .Y(_00747_));
 sky130_fd_sc_hd__nand3_1 _06931_ (.A(_00576_),
    .B(net44),
    .C(net14),
    .Y(_00749_));
 sky130_fd_sc_hd__o2111ai_4 _06932_ (.A1(_00414_),
    .A2(_00744_),
    .B1(net13),
    .C1(net55),
    .D1(_00746_),
    .Y(_00750_));
 sky130_fd_sc_hd__o21ai_2 _06933_ (.A1(_00414_),
    .A2(_00744_),
    .B1(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__a21oi_1 _06934_ (.A1(_00577_),
    .A2(_00581_),
    .B1(_00578_),
    .Y(_00752_));
 sky130_fd_sc_hd__o2bb2ai_2 _06935_ (.A1_N(_00577_),
    .A2_N(_00581_),
    .B1(_00242_),
    .B2(_00341_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(_00751_),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand3_4 _06937_ (.A(_00584_),
    .B(_00751_),
    .C(_00753_),
    .Y(_00755_));
 sky130_fd_sc_hd__a21oi_1 _06938_ (.A1(_00584_),
    .A2(_00753_),
    .B1(_00751_),
    .Y(_00756_));
 sky130_fd_sc_hd__o21bai_4 _06939_ (.A1(_00582_),
    .A2(_00752_),
    .B1_N(_00751_),
    .Y(_00757_));
 sky130_fd_sc_hd__a22o_1 _06940_ (.A1(net13),
    .A2(net58),
    .B1(net59),
    .B2(net11),
    .X(_00758_));
 sky130_fd_sc_hd__and3_1 _06941_ (.A(net11),
    .B(net13),
    .C(net58),
    .X(_00760_));
 sky130_fd_sc_hd__and4_1 _06942_ (.A(net11),
    .B(net13),
    .C(net58),
    .D(net59),
    .X(_00761_));
 sky130_fd_sc_hd__a21bo_1 _06943_ (.A1(net59),
    .A2(_00760_),
    .B1_N(_00758_),
    .X(_00762_));
 sky130_fd_sc_hd__and4b_1 _06944_ (.A_N(_00761_),
    .B(net60),
    .C(net10),
    .D(_00758_),
    .X(_00763_));
 sky130_fd_sc_hd__o21a_1 _06945_ (.A1(_00231_),
    .A2(_00352_),
    .B1(_00762_),
    .X(_00764_));
 sky130_fd_sc_hd__a21oi_2 _06946_ (.A1(net10),
    .A2(net60),
    .B1(_00762_),
    .Y(_00765_));
 sky130_fd_sc_hd__and3_1 _06947_ (.A(_00762_),
    .B(net60),
    .C(net10),
    .X(_00766_));
 sky130_fd_sc_hd__nor2_1 _06948_ (.A(_00765_),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__o211ai_4 _06949_ (.A1(_00765_),
    .A2(_00766_),
    .B1(_00755_),
    .C1(_00757_),
    .Y(_00768_));
 sky130_fd_sc_hd__o22ai_4 _06950_ (.A1(_00582_),
    .A2(_00754_),
    .B1(_00767_),
    .B2(_00756_),
    .Y(_00769_));
 sky130_fd_sc_hd__o2bb2ai_1 _06951_ (.A1_N(_00587_),
    .A2_N(_00588_),
    .B1(_00595_),
    .B2(_00596_),
    .Y(_00771_));
 sky130_fd_sc_hd__o211ai_2 _06952_ (.A1(_00592_),
    .A2(_00593_),
    .B1(_00587_),
    .C1(_00588_),
    .Y(_00772_));
 sky130_fd_sc_hd__o221a_1 _06953_ (.A1(_00574_),
    .A2(_00585_),
    .B1(_00595_),
    .B2(_00596_),
    .C1(_00587_),
    .X(_00773_));
 sky130_fd_sc_hd__o221ai_4 _06954_ (.A1(_00574_),
    .A2(_00585_),
    .B1(_00595_),
    .B2(_00596_),
    .C1(_00587_),
    .Y(_00774_));
 sky130_fd_sc_hd__o2bb2ai_4 _06955_ (.A1_N(_00587_),
    .A2_N(_00588_),
    .B1(_00592_),
    .B2(_00593_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(_00769_),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand3_4 _06957_ (.A(_00769_),
    .B(_00774_),
    .C(_00775_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _06958_ (.A(net8),
    .B(net61),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _06959_ (.A(net8),
    .B(net62),
    .Y(_00779_));
 sky130_fd_sc_hd__and4_1 _06960_ (.A(net9),
    .B(net8),
    .C(net62),
    .D(net61),
    .X(_00780_));
 sky130_fd_sc_hd__a22o_1 _06961_ (.A1(net8),
    .A2(net62),
    .B1(net61),
    .B2(net9),
    .X(_00782_));
 sky130_fd_sc_hd__nand3_1 _06962_ (.A(_00779_),
    .B(net61),
    .C(net9),
    .Y(_00783_));
 sky130_fd_sc_hd__nand3_1 _06963_ (.A(_00601_),
    .B(net62),
    .C(net8),
    .Y(_00784_));
 sky130_fd_sc_hd__o2111ai_2 _06964_ (.A1(_00602_),
    .A2(_00778_),
    .B1(net7),
    .C1(net63),
    .D1(_00782_),
    .Y(_00785_));
 sky130_fd_sc_hd__a31o_1 _06965_ (.A1(_00782_),
    .A2(net63),
    .A3(net7),
    .B1(_00780_),
    .X(_00786_));
 sky130_fd_sc_hd__a31o_1 _06966_ (.A1(_00758_),
    .A2(net60),
    .A3(net10),
    .B1(_00761_),
    .X(_00787_));
 sky130_fd_sc_hd__o22ai_2 _06967_ (.A1(_00209_),
    .A2(_00396_),
    .B1(_00603_),
    .B2(_00604_),
    .Y(_00788_));
 sky130_fd_sc_hd__a21o_1 _06968_ (.A1(_00608_),
    .A2(_00788_),
    .B1(_00787_),
    .X(_00789_));
 sky130_fd_sc_hd__nand3_4 _06969_ (.A(_00608_),
    .B(_00787_),
    .C(_00788_),
    .Y(_00790_));
 sky130_fd_sc_hd__and2_1 _06970_ (.A(_00789_),
    .B(_00790_),
    .X(_00791_));
 sky130_fd_sc_hd__nand3_4 _06971_ (.A(_00786_),
    .B(_00789_),
    .C(_00790_),
    .Y(_00793_));
 sky130_fd_sc_hd__a311o_1 _06972_ (.A1(net7),
    .A2(_00782_),
    .A3(net63),
    .B1(_00780_),
    .C1(_00791_),
    .X(_00794_));
 sky130_fd_sc_hd__a21boi_2 _06973_ (.A1(_00789_),
    .A2(_00790_),
    .B1_N(_00786_),
    .Y(_00795_));
 sky130_fd_sc_hd__o311a_1 _06974_ (.A1(_00209_),
    .A2(_00385_),
    .A3(_00602_),
    .B1(_00785_),
    .C1(_00791_),
    .X(_00796_));
 sky130_fd_sc_hd__nor2_1 _06975_ (.A(_00795_),
    .B(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__a21oi_4 _06976_ (.A1(_00774_),
    .A2(_00775_),
    .B1(_00769_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand4_4 _06977_ (.A(_00755_),
    .B(_00768_),
    .C(_00771_),
    .D(_00772_),
    .Y(_00799_));
 sky130_fd_sc_hd__o21ai_1 _06978_ (.A1(_00795_),
    .A2(_00796_),
    .B1(_00777_),
    .Y(_00800_));
 sky130_fd_sc_hd__o211a_4 _06979_ (.A1(_00795_),
    .A2(_00796_),
    .B1(_00799_),
    .C1(_00777_),
    .X(_00801_));
 sky130_fd_sc_hd__o22a_1 _06980_ (.A1(_00773_),
    .A2(_00776_),
    .B1(_00797_),
    .B2(_00798_),
    .X(_00802_));
 sky130_fd_sc_hd__o21ai_1 _06981_ (.A1(_00797_),
    .A2(_00798_),
    .B1(_00777_),
    .Y(_00804_));
 sky130_fd_sc_hd__a21o_1 _06982_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_00618_),
    .X(_00805_));
 sky130_fd_sc_hd__o211a_1 _06983_ (.A1(_00614_),
    .A2(_00617_),
    .B1(_00599_),
    .C1(_00600_),
    .X(_00806_));
 sky130_fd_sc_hd__a211oi_2 _06984_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_00614_),
    .C1(_00617_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(_00619_),
    .B(_00805_),
    .Y(_00808_));
 sky130_fd_sc_hd__a32o_2 _06986_ (.A1(_00769_),
    .A2(_00774_),
    .A3(_00775_),
    .B1(_00805_),
    .B2(_00619_),
    .X(_00809_));
 sky130_fd_sc_hd__o211ai_4 _06987_ (.A1(_00798_),
    .A2(_00797_),
    .B1(_00777_),
    .C1(_00808_),
    .Y(_00810_));
 sky130_fd_sc_hd__o21ai_4 _06988_ (.A1(_00806_),
    .A2(_00807_),
    .B1(_00804_),
    .Y(_00811_));
 sky130_fd_sc_hd__a22o_1 _06989_ (.A1(net5),
    .A2(net35),
    .B1(_00626_),
    .B2(_00628_),
    .X(_00812_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(net5),
    .B(net64),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(net5),
    .B(net34),
    .Y(_00815_));
 sky130_fd_sc_hd__and4_1 _06992_ (.A(net5),
    .B(net6),
    .C(net64),
    .D(net34),
    .X(_00816_));
 sky130_fd_sc_hd__nand4_2 _06993_ (.A(net5),
    .B(net6),
    .C(net64),
    .D(net34),
    .Y(_00817_));
 sky130_fd_sc_hd__a22oi_4 _06994_ (.A1(net6),
    .A2(net64),
    .B1(net34),
    .B2(net5),
    .Y(_00818_));
 sky130_fd_sc_hd__nand4b_2 _06995_ (.A_N(_00818_),
    .B(net35),
    .C(net4),
    .D(_00817_),
    .Y(_00819_));
 sky130_fd_sc_hd__o31ai_4 _06996_ (.A1(_00165_),
    .A2(_00407_),
    .A3(_00818_),
    .B1(_00817_),
    .Y(_00820_));
 sky130_fd_sc_hd__o211a_1 _06997_ (.A1(_00154_),
    .A2(_00630_),
    .B1(_00812_),
    .C1(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__o211ai_4 _06998_ (.A1(_00154_),
    .A2(_00630_),
    .B1(_00812_),
    .C1(_00820_),
    .Y(_00822_));
 sky130_fd_sc_hd__a22oi_2 _06999_ (.A1(net2),
    .A2(net38),
    .B1(_00665_),
    .B2(_00667_),
    .Y(_00823_));
 sky130_fd_sc_hd__nor2_1 _07000_ (.A(_00669_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__a21oi_1 _07001_ (.A1(_00631_),
    .A2(_00812_),
    .B1(_00820_),
    .Y(_00826_));
 sky130_fd_sc_hd__a21o_1 _07002_ (.A1(_00631_),
    .A2(_00812_),
    .B1(_00820_),
    .X(_00827_));
 sky130_fd_sc_hd__or3b_2 _07003_ (.A(_00821_),
    .B(_00826_),
    .C_N(_00824_),
    .X(_00828_));
 sky130_fd_sc_hd__o31a_1 _07004_ (.A1(_00669_),
    .A2(_00823_),
    .A3(_00826_),
    .B1(_00822_),
    .X(_00829_));
 sky130_fd_sc_hd__a21o_1 _07005_ (.A1(_00827_),
    .A2(_00824_),
    .B1(_00821_),
    .X(_00830_));
 sky130_fd_sc_hd__a21bo_1 _07006_ (.A1(_00786_),
    .A2(_00789_),
    .B1_N(_00790_),
    .X(_00831_));
 sky130_fd_sc_hd__a22oi_4 _07007_ (.A1(_00502_),
    .A2(_00636_),
    .B1(_00640_),
    .B2(_00635_),
    .Y(_00832_));
 sky130_fd_sc_hd__o2bb2ai_1 _07008_ (.A1_N(_00502_),
    .A2_N(_00636_),
    .B1(_00639_),
    .B2(_00634_),
    .Y(_00833_));
 sky130_fd_sc_hd__a211oi_4 _07009_ (.A1(_00790_),
    .A2(_00793_),
    .B1(_00832_),
    .C1(_00641_),
    .Y(_00834_));
 sky130_fd_sc_hd__a211o_1 _07010_ (.A1(_00790_),
    .A2(_00793_),
    .B1(_00832_),
    .C1(_00641_),
    .X(_00835_));
 sky130_fd_sc_hd__a21oi_2 _07011_ (.A1(_00642_),
    .A2(_00833_),
    .B1(_00831_),
    .Y(_00837_));
 sky130_fd_sc_hd__a211oi_4 _07012_ (.A1(_00822_),
    .A2(_00828_),
    .B1(_00834_),
    .C1(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__o211a_2 _07013_ (.A1(_00834_),
    .A2(_00837_),
    .B1(_00822_),
    .C1(_00828_),
    .X(_00839_));
 sky130_fd_sc_hd__o2bb2a_1 _07014_ (.A1_N(_00822_),
    .A2_N(_00828_),
    .B1(_00834_),
    .B2(_00837_),
    .X(_00840_));
 sky130_fd_sc_hd__or3_1 _07015_ (.A(_00830_),
    .B(_00834_),
    .C(_00837_),
    .X(_00841_));
 sky130_fd_sc_hd__inv_2 _07016_ (.A(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _07017_ (.A(_00838_),
    .B(_00839_),
    .Y(_00843_));
 sky130_fd_sc_hd__o22ai_2 _07018_ (.A1(_00838_),
    .A2(_00839_),
    .B1(_00808_),
    .B2(_00802_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_00810_),
    .B(_00843_),
    .Y(_00845_));
 sky130_fd_sc_hd__o2111ai_4 _07020_ (.A1(_00801_),
    .A2(_00809_),
    .B1(_00844_),
    .C1(_00741_),
    .D1(_00658_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand4_2 _07021_ (.A(_00742_),
    .B(_00743_),
    .C(_00811_),
    .D(_00845_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand4_1 _07022_ (.A(_00658_),
    .B(_00741_),
    .C(_00811_),
    .D(_00845_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand4_1 _07023_ (.A(_00742_),
    .B(_00743_),
    .C(_00810_),
    .D(_00844_),
    .Y(_00850_));
 sky130_fd_sc_hd__o22ai_4 _07024_ (.A1(_00088_),
    .A2(_00451_),
    .B1(_00676_),
    .B2(_00677_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _07025_ (.A(net2),
    .B(net36),
    .Y(_00852_));
 sky130_fd_sc_hd__or2_1 _07026_ (.A(_00666_),
    .B(_00852_),
    .X(_00853_));
 sky130_fd_sc_hd__and2_1 _07027_ (.A(net32),
    .B(net38),
    .X(_00854_));
 sky130_fd_sc_hd__a22o_1 _07028_ (.A1(net2),
    .A2(net37),
    .B1(net36),
    .B2(net3),
    .X(_00855_));
 sky130_fd_sc_hd__o311a_1 _07029_ (.A1(_00143_),
    .A2(_00429_),
    .A3(_00666_),
    .B1(_00854_),
    .C1(_00855_),
    .X(_00856_));
 sky130_fd_sc_hd__o2bb2ai_2 _07030_ (.A1_N(_00854_),
    .A2_N(_00855_),
    .B1(_00666_),
    .B2(_00852_),
    .Y(_00857_));
 sky130_fd_sc_hd__and3_1 _07031_ (.A(_00679_),
    .B(_00851_),
    .C(_00857_),
    .X(_00859_));
 sky130_fd_sc_hd__nand3_2 _07032_ (.A(_00679_),
    .B(_00851_),
    .C(_00857_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand2_2 _07033_ (.A(net30),
    .B(net40),
    .Y(_00861_));
 sky130_fd_sc_hd__nand4_2 _07034_ (.A(net30),
    .B(net31),
    .C(net39),
    .D(net40),
    .Y(_00862_));
 sky130_fd_sc_hd__a22o_1 _07035_ (.A1(net31),
    .A2(net39),
    .B1(net40),
    .B2(net30),
    .X(_00863_));
 sky130_fd_sc_hd__nand3_1 _07036_ (.A(_00861_),
    .B(net39),
    .C(net31),
    .Y(_00864_));
 sky130_fd_sc_hd__nand3_1 _07037_ (.A(_00675_),
    .B(net40),
    .C(net30),
    .Y(_00865_));
 sky130_fd_sc_hd__nand4_4 _07038_ (.A(_00863_),
    .B(net41),
    .C(net29),
    .D(_00862_),
    .Y(_00866_));
 sky130_fd_sc_hd__o31a_1 _07039_ (.A1(_00121_),
    .A2(_00440_),
    .A3(_00861_),
    .B1(_00866_),
    .X(_00867_));
 sky130_fd_sc_hd__o21ai_1 _07040_ (.A1(_00675_),
    .A2(_00861_),
    .B1(_00866_),
    .Y(_00868_));
 sky130_fd_sc_hd__a21oi_2 _07041_ (.A1(_00679_),
    .A2(_00851_),
    .B1(_00857_),
    .Y(_00870_));
 sky130_fd_sc_hd__a21o_1 _07042_ (.A1(_00679_),
    .A2(_00851_),
    .B1(_00857_),
    .X(_00871_));
 sky130_fd_sc_hd__o21a_1 _07043_ (.A1(_00867_),
    .A2(_00870_),
    .B1(_00860_),
    .X(_00872_));
 sky130_fd_sc_hd__o21ai_1 _07044_ (.A1(_00867_),
    .A2(_00870_),
    .B1(_00860_),
    .Y(_00873_));
 sky130_fd_sc_hd__o21bai_1 _07045_ (.A1(_00673_),
    .A2(_00681_),
    .B1_N(_00680_),
    .Y(_00874_));
 sky130_fd_sc_hd__o21ai_1 _07046_ (.A1(_00673_),
    .A2(_00681_),
    .B1(_00680_),
    .Y(_00875_));
 sky130_fd_sc_hd__nand3b_1 _07047_ (.A_N(_00680_),
    .B(_00683_),
    .C(_00674_),
    .Y(_00876_));
 sky130_fd_sc_hd__and3_1 _07048_ (.A(_00684_),
    .B(_00873_),
    .C(_00874_),
    .X(_00877_));
 sky130_fd_sc_hd__nand3_1 _07049_ (.A(_00684_),
    .B(_00873_),
    .C(_00874_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand3_1 _07050_ (.A(_00872_),
    .B(_00875_),
    .C(_00876_),
    .Y(_00879_));
 sky130_fd_sc_hd__a22oi_1 _07051_ (.A1(net27),
    .A2(net46),
    .B1(net47),
    .B2(net26),
    .Y(_00881_));
 sky130_fd_sc_hd__a22o_1 _07052_ (.A1(net27),
    .A2(net46),
    .B1(net47),
    .B2(net26),
    .X(_00882_));
 sky130_fd_sc_hd__nand4_2 _07053_ (.A(net26),
    .B(net27),
    .C(net46),
    .D(net47),
    .Y(_00883_));
 sky130_fd_sc_hd__a22o_1 _07054_ (.A1(_00882_),
    .A2(_00883_),
    .B1(net117),
    .B2(net23),
    .X(_00884_));
 sky130_fd_sc_hd__nand4b_2 _07055_ (.A_N(_00881_),
    .B(net23),
    .C(net117),
    .D(_00883_),
    .Y(_00885_));
 sky130_fd_sc_hd__and4_1 _07056_ (.A(net28),
    .B(net29),
    .C(net43),
    .D(net42),
    .X(_00886_));
 sky130_fd_sc_hd__nand4_1 _07057_ (.A(net28),
    .B(net29),
    .C(net43),
    .D(net42),
    .Y(_00887_));
 sky130_fd_sc_hd__a22o_1 _07058_ (.A1(net28),
    .A2(net43),
    .B1(net42),
    .B2(net29),
    .X(_00888_));
 sky130_fd_sc_hd__nand4_2 _07059_ (.A(_00888_),
    .B(net45),
    .C(net27),
    .D(_00887_),
    .Y(_00889_));
 sky130_fd_sc_hd__a31o_1 _07060_ (.A1(_00888_),
    .A2(net45),
    .A3(net27),
    .B1(_00886_),
    .X(_00890_));
 sky130_fd_sc_hd__a22o_1 _07061_ (.A1(net28),
    .A2(net45),
    .B1(_00695_),
    .B2(_00696_),
    .X(_00892_));
 sky130_fd_sc_hd__a21o_1 _07062_ (.A1(_00697_),
    .A2(_00892_),
    .B1(_00890_),
    .X(_00893_));
 sky130_fd_sc_hd__and3_1 _07063_ (.A(_00697_),
    .B(_00890_),
    .C(_00892_),
    .X(_00894_));
 sky130_fd_sc_hd__nand3_1 _07064_ (.A(_00697_),
    .B(_00890_),
    .C(_00892_),
    .Y(_00895_));
 sky130_fd_sc_hd__and4_1 _07065_ (.A(_00884_),
    .B(_00885_),
    .C(_00893_),
    .D(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__nand4_1 _07066_ (.A(_00884_),
    .B(_00885_),
    .C(_00893_),
    .D(_00895_),
    .Y(_00897_));
 sky130_fd_sc_hd__a22o_1 _07067_ (.A1(_00884_),
    .A2(_00885_),
    .B1(_00893_),
    .B2(_00895_),
    .X(_00898_));
 sky130_fd_sc_hd__nand2_1 _07068_ (.A(_00897_),
    .B(_00898_),
    .Y(_00899_));
 sky130_fd_sc_hd__a31o_1 _07069_ (.A1(_00879_),
    .A2(_00897_),
    .A3(_00898_),
    .B1(_00877_),
    .X(_00900_));
 sky130_fd_sc_hd__inv_2 _07070_ (.A(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__o21ai_1 _07071_ (.A1(_00829_),
    .A2(_00837_),
    .B1(_00835_),
    .Y(_00903_));
 sky130_fd_sc_hd__a22o_1 _07072_ (.A1(_00701_),
    .A2(_00702_),
    .B1(_00705_),
    .B2(_00688_),
    .X(_00904_));
 sky130_fd_sc_hd__a21o_1 _07073_ (.A1(_00688_),
    .A2(_00705_),
    .B1(_00703_),
    .X(_00905_));
 sky130_fd_sc_hd__nand3_1 _07074_ (.A(_00688_),
    .B(_00703_),
    .C(_00705_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand3_1 _07075_ (.A(_00706_),
    .B(_00903_),
    .C(_00904_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand3b_1 _07076_ (.A_N(_00903_),
    .B(_00905_),
    .C(_00906_),
    .Y(_00908_));
 sky130_fd_sc_hd__a21oi_1 _07077_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00901_),
    .Y(_00909_));
 sky130_fd_sc_hd__and3_1 _07078_ (.A(_00901_),
    .B(_00907_),
    .C(_00908_),
    .X(_00910_));
 sky130_fd_sc_hd__nor2_1 _07079_ (.A(_00909_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__o211ai_2 _07080_ (.A1(_00909_),
    .A2(_00910_),
    .B1(_00846_),
    .C1(_00848_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _07081_ (.A(_00846_),
    .B(_00912_),
    .Y(_00914_));
 sky130_fd_sc_hd__a22o_1 _07082_ (.A1(_00663_),
    .A2(_00664_),
    .B1(_00712_),
    .B2(_00713_),
    .X(_00915_));
 sky130_fd_sc_hd__a21oi_1 _07083_ (.A1(_00714_),
    .A2(_00915_),
    .B1(_00914_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _07084_ (.A(_00714_),
    .B(_00914_),
    .C(_00915_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _07085_ (.A(_00690_),
    .B(_00692_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_1 _07086_ (.A(_00700_),
    .B(_00702_),
    .Y(_00919_));
 sky130_fd_sc_hd__a21bo_1 _07087_ (.A1(_00900_),
    .A2(_00908_),
    .B1_N(_00907_),
    .X(_00920_));
 sky130_fd_sc_hd__xor2_1 _07088_ (.A(_00919_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__xnor2_1 _07089_ (.A(_00918_),
    .B(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__or2_1 _07090_ (.A(_00916_),
    .B(_00922_),
    .X(_00923_));
 sky130_fd_sc_hd__nor3_1 _07091_ (.A(_00717_),
    .B(_00718_),
    .C(_00725_),
    .Y(_00925_));
 sky130_fd_sc_hd__o21a_1 _07092_ (.A1(_00717_),
    .A2(_00718_),
    .B1(_00725_),
    .X(_00926_));
 sky130_fd_sc_hd__a211o_1 _07093_ (.A1(_00917_),
    .A2(_00923_),
    .B1(_00925_),
    .C1(_00926_),
    .X(_00927_));
 sky130_fd_sc_hd__a22oi_2 _07094_ (.A1(_00919_),
    .A2(_00920_),
    .B1(_00921_),
    .B2(_00918_),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _07095_ (.A(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__o221a_1 _07096_ (.A1(_00916_),
    .A2(_00922_),
    .B1(_00925_),
    .B2(_00926_),
    .C1(_00917_),
    .X(_00930_));
 sky130_fd_sc_hd__inv_2 _07097_ (.A(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _07098_ (.A(_00927_),
    .B(_00929_),
    .Y(_00932_));
 sky130_fd_sc_hd__and3_1 _07099_ (.A(_00927_),
    .B(_00929_),
    .C(_00931_),
    .X(_00933_));
 sky130_fd_sc_hd__o21a_1 _07100_ (.A1(_00928_),
    .A2(_00930_),
    .B1(_00927_),
    .X(_00934_));
 sky130_fd_sc_hd__nand2_1 _07101_ (.A(_00731_),
    .B(_00729_),
    .Y(_00936_));
 sky130_fd_sc_hd__o21ba_1 _07102_ (.A1(_00729_),
    .A2(_00731_),
    .B1_N(_00934_),
    .X(_00937_));
 sky130_fd_sc_hd__a21oi_1 _07103_ (.A1(_00927_),
    .A2(_00931_),
    .B1(_00929_),
    .Y(_00938_));
 sky130_fd_sc_hd__o21bai_1 _07104_ (.A1(_00930_),
    .A2(_00932_),
    .B1_N(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__o2bb2ai_4 _07105_ (.A1_N(_00755_),
    .A2_N(_00757_),
    .B1(_00763_),
    .B2(_00764_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_2 _07106_ (.A(net13),
    .B(net33),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_2 _07107_ (.A(net13),
    .B(net44),
    .Y(_00942_));
 sky130_fd_sc_hd__and4_1 _07108_ (.A(net14),
    .B(net13),
    .C(net44),
    .D(net33),
    .X(_00943_));
 sky130_fd_sc_hd__nand2_1 _07109_ (.A(net11),
    .B(net55),
    .Y(_00944_));
 sky130_fd_sc_hd__a22oi_2 _07110_ (.A1(net13),
    .A2(net44),
    .B1(net33),
    .B2(net14),
    .Y(_00945_));
 sky130_fd_sc_hd__a22o_1 _07111_ (.A1(net13),
    .A2(net44),
    .B1(net33),
    .B2(net14),
    .X(_00947_));
 sky130_fd_sc_hd__nand3_1 _07112_ (.A(_00942_),
    .B(net33),
    .C(net14),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3_1 _07113_ (.A(_00744_),
    .B(net44),
    .C(net13),
    .Y(_00949_));
 sky130_fd_sc_hd__o2111ai_4 _07114_ (.A1(_00745_),
    .A2(_00941_),
    .B1(net11),
    .C1(net55),
    .D1(_00947_),
    .Y(_00950_));
 sky130_fd_sc_hd__o22ai_2 _07115_ (.A1(_00745_),
    .A2(_00941_),
    .B1(_00944_),
    .B2(_00945_),
    .Y(_00951_));
 sky130_fd_sc_hd__o211ai_2 _07116_ (.A1(_00253_),
    .A2(_00341_),
    .B1(_00747_),
    .C1(_00749_),
    .Y(_00952_));
 sky130_fd_sc_hd__and3_1 _07117_ (.A(_00750_),
    .B(_00951_),
    .C(_00952_),
    .X(_00953_));
 sky130_fd_sc_hd__nand3_2 _07118_ (.A(_00750_),
    .B(_00951_),
    .C(_00952_),
    .Y(_00954_));
 sky130_fd_sc_hd__a21o_2 _07119_ (.A1(_00750_),
    .A2(_00952_),
    .B1(_00951_),
    .X(_00955_));
 sky130_fd_sc_hd__inv_2 _07120_ (.A(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__and4_1 _07121_ (.A(net11),
    .B(net10),
    .C(net58),
    .D(net59),
    .X(_00958_));
 sky130_fd_sc_hd__nand4_1 _07122_ (.A(net11),
    .B(net10),
    .C(net58),
    .D(net59),
    .Y(_00959_));
 sky130_fd_sc_hd__a22oi_4 _07123_ (.A1(net11),
    .A2(net58),
    .B1(net59),
    .B2(net10),
    .Y(_00960_));
 sky130_fd_sc_hd__and4b_1 _07124_ (.A_N(_00960_),
    .B(net60),
    .C(net9),
    .D(_00959_),
    .X(_00961_));
 sky130_fd_sc_hd__o22a_1 _07125_ (.A1(_00198_),
    .A2(_00352_),
    .B1(_00958_),
    .B2(_00960_),
    .X(_00962_));
 sky130_fd_sc_hd__a211oi_2 _07126_ (.A1(net9),
    .A2(net60),
    .B1(_00958_),
    .C1(_00960_),
    .Y(_00963_));
 sky130_fd_sc_hd__a211o_1 _07127_ (.A1(net9),
    .A2(net60),
    .B1(_00958_),
    .C1(_00960_),
    .X(_00964_));
 sky130_fd_sc_hd__o211a_1 _07128_ (.A1(_00958_),
    .A2(_00960_),
    .B1(net9),
    .C1(net60),
    .X(_00965_));
 sky130_fd_sc_hd__o211ai_1 _07129_ (.A1(_00958_),
    .A2(_00960_),
    .B1(net9),
    .C1(net60),
    .Y(_00966_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(_00964_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__and3_1 _07131_ (.A(_00954_),
    .B(_00964_),
    .C(_00966_),
    .X(_00969_));
 sky130_fd_sc_hd__o31a_1 _07132_ (.A1(_00953_),
    .A2(_00963_),
    .A3(_00965_),
    .B1(_00955_),
    .X(_00970_));
 sky130_fd_sc_hd__a21oi_2 _07133_ (.A1(_00768_),
    .A2(_00940_),
    .B1(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__o2bb2ai_4 _07134_ (.A1_N(_00768_),
    .A2_N(_00940_),
    .B1(_00956_),
    .B2(_00969_),
    .Y(_00972_));
 sky130_fd_sc_hd__o2111ai_4 _07135_ (.A1(_00953_),
    .A2(_00967_),
    .B1(_00955_),
    .C1(_00768_),
    .D1(_00940_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand4_4 _07136_ (.A(net7),
    .B(net8),
    .C(net62),
    .D(net61),
    .Y(_00974_));
 sky130_fd_sc_hd__a22o_1 _07137_ (.A1(net7),
    .A2(net62),
    .B1(net61),
    .B2(net8),
    .X(_00975_));
 sky130_fd_sc_hd__nand4_4 _07138_ (.A(_00975_),
    .B(net63),
    .C(net6),
    .D(_00974_),
    .Y(_00976_));
 sky130_fd_sc_hd__o31a_1 _07139_ (.A1(_00176_),
    .A2(_00374_),
    .A3(_00778_),
    .B1(_00976_),
    .X(_00977_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(_00974_),
    .B(_00976_),
    .Y(_00978_));
 sky130_fd_sc_hd__o31ai_2 _07141_ (.A1(_00198_),
    .A2(_00352_),
    .A3(_00960_),
    .B1(_00959_),
    .Y(_00980_));
 sky130_fd_sc_hd__o211ai_1 _07142_ (.A1(_00176_),
    .A2(_00396_),
    .B1(_00783_),
    .C1(_00784_),
    .Y(_00981_));
 sky130_fd_sc_hd__a21oi_1 _07143_ (.A1(_00785_),
    .A2(_00981_),
    .B1(_00980_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand3_1 _07144_ (.A(_00785_),
    .B(_00980_),
    .C(_00981_),
    .Y(_00983_));
 sky130_fd_sc_hd__and2b_1 _07145_ (.A_N(_00982_),
    .B(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__and2_1 _07146_ (.A(_00984_),
    .B(_00978_),
    .X(_00985_));
 sky130_fd_sc_hd__nor2_2 _07147_ (.A(_00978_),
    .B(_00984_),
    .Y(_00986_));
 sky130_fd_sc_hd__a21oi_1 _07148_ (.A1(_00974_),
    .A2(_00976_),
    .B1(_00984_),
    .Y(_00987_));
 sky130_fd_sc_hd__o311a_1 _07149_ (.A1(_00176_),
    .A2(_00385_),
    .A3(_00779_),
    .B1(_00976_),
    .C1(_00984_),
    .X(_00988_));
 sky130_fd_sc_hd__nor2_1 _07150_ (.A(_00985_),
    .B(_00986_),
    .Y(_00989_));
 sky130_fd_sc_hd__a31oi_2 _07151_ (.A1(_00768_),
    .A2(_00940_),
    .A3(_00970_),
    .B1(_00989_),
    .Y(_00991_));
 sky130_fd_sc_hd__a31o_1 _07152_ (.A1(_00768_),
    .A2(_00940_),
    .A3(_00970_),
    .B1(_00989_),
    .X(_00992_));
 sky130_fd_sc_hd__a22oi_4 _07153_ (.A1(_00793_),
    .A2(_00794_),
    .B1(_00799_),
    .B2(_00777_),
    .Y(_00993_));
 sky130_fd_sc_hd__a22o_1 _07154_ (.A1(_00793_),
    .A2(_00794_),
    .B1(_00799_),
    .B2(_00777_),
    .X(_00994_));
 sky130_fd_sc_hd__o22a_1 _07155_ (.A1(_00971_),
    .A2(_00991_),
    .B1(_00993_),
    .B2(_00801_),
    .X(_00995_));
 sky130_fd_sc_hd__o22ai_4 _07156_ (.A1(_00971_),
    .A2(_00991_),
    .B1(_00993_),
    .B2(_00801_),
    .Y(_00996_));
 sky130_fd_sc_hd__o2111ai_4 _07157_ (.A1(_00798_),
    .A2(_00800_),
    .B1(_00972_),
    .C1(_00992_),
    .D1(_00994_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _07158_ (.A(net4),
    .B(net64),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(net4),
    .B(net34),
    .Y(_00999_));
 sky130_fd_sc_hd__and2_1 _07160_ (.A(net3),
    .B(net35),
    .X(_01000_));
 sky130_fd_sc_hd__a22o_1 _07161_ (.A1(net5),
    .A2(net64),
    .B1(net34),
    .B2(net4),
    .X(_01002_));
 sky130_fd_sc_hd__nand3_1 _07162_ (.A(_00999_),
    .B(net64),
    .C(net5),
    .Y(_01003_));
 sky130_fd_sc_hd__nand3_1 _07163_ (.A(_00813_),
    .B(net34),
    .C(net4),
    .Y(_01004_));
 sky130_fd_sc_hd__o2111ai_4 _07164_ (.A1(_00815_),
    .A2(_00998_),
    .B1(net3),
    .C1(net35),
    .D1(_01002_),
    .Y(_01005_));
 sky130_fd_sc_hd__o2bb2ai_2 _07165_ (.A1_N(_01000_),
    .A2_N(_01002_),
    .B1(_00815_),
    .B2(_00998_),
    .Y(_01006_));
 sky130_fd_sc_hd__o22a_1 _07166_ (.A1(_00165_),
    .A2(_00407_),
    .B1(_00816_),
    .B2(_00818_),
    .X(_01007_));
 sky130_fd_sc_hd__o22ai_2 _07167_ (.A1(_00165_),
    .A2(_00407_),
    .B1(_00816_),
    .B2(_00818_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(_00819_),
    .B(_01006_),
    .Y(_01009_));
 sky130_fd_sc_hd__and3_1 _07169_ (.A(_00819_),
    .B(_01006_),
    .C(_01008_),
    .X(_01010_));
 sky130_fd_sc_hd__a21oi_1 _07170_ (.A1(_00853_),
    .A2(_00855_),
    .B1(_00854_),
    .Y(_01011_));
 sky130_fd_sc_hd__nor2_1 _07171_ (.A(_00856_),
    .B(_01011_),
    .Y(_01013_));
 sky130_fd_sc_hd__a21oi_1 _07172_ (.A1(_00819_),
    .A2(_01008_),
    .B1(_01006_),
    .Y(_01014_));
 sky130_fd_sc_hd__a21o_1 _07173_ (.A1(_00819_),
    .A2(_01008_),
    .B1(_01006_),
    .X(_01015_));
 sky130_fd_sc_hd__o211ai_2 _07174_ (.A1(_01007_),
    .A2(_01009_),
    .B1(_01015_),
    .C1(_01013_),
    .Y(_01016_));
 sky130_fd_sc_hd__o32a_1 _07175_ (.A1(_00856_),
    .A2(_01011_),
    .A3(_01014_),
    .B1(_01007_),
    .B2(_01009_),
    .X(_01017_));
 sky130_fd_sc_hd__a2bb2o_1 _07176_ (.A1_N(_01007_),
    .A2_N(_01009_),
    .B1(_01015_),
    .B2(_01013_),
    .X(_01018_));
 sky130_fd_sc_hd__o21ai_2 _07177_ (.A1(_00977_),
    .A2(_00982_),
    .B1(_00983_),
    .Y(_01019_));
 sky130_fd_sc_hd__o21ai_2 _07178_ (.A1(_00821_),
    .A2(_00826_),
    .B1(_00824_),
    .Y(_01020_));
 sky130_fd_sc_hd__o211ai_2 _07179_ (.A1(_00669_),
    .A2(_00823_),
    .B1(_00827_),
    .C1(_00822_),
    .Y(_01021_));
 sky130_fd_sc_hd__a21boi_1 _07180_ (.A1(_01020_),
    .A2(_01021_),
    .B1_N(_01019_),
    .Y(_01022_));
 sky130_fd_sc_hd__a21bo_1 _07181_ (.A1(_01020_),
    .A2(_01021_),
    .B1_N(_01019_),
    .X(_01024_));
 sky130_fd_sc_hd__nand3b_2 _07182_ (.A_N(_01019_),
    .B(_01020_),
    .C(_01021_),
    .Y(_01025_));
 sky130_fd_sc_hd__and3_2 _07183_ (.A(_01018_),
    .B(_01024_),
    .C(_01025_),
    .X(_01026_));
 sky130_fd_sc_hd__a21oi_2 _07184_ (.A1(_01024_),
    .A2(_01025_),
    .B1(_01018_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21oi_2 _07185_ (.A1(_01024_),
    .A2(_01025_),
    .B1(_01017_),
    .Y(_01028_));
 sky130_fd_sc_hd__and3_1 _07186_ (.A(_01024_),
    .B(_01025_),
    .C(_01017_),
    .X(_01029_));
 sky130_fd_sc_hd__nor2_1 _07187_ (.A(_01028_),
    .B(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__o21ai_2 _07188_ (.A1(_01026_),
    .A2(_01027_),
    .B1(_00997_),
    .Y(_01031_));
 sky130_fd_sc_hd__o221ai_4 _07189_ (.A1(_00838_),
    .A2(_00839_),
    .B1(_00801_),
    .B2(_00809_),
    .C1(_00811_),
    .Y(_01032_));
 sky130_fd_sc_hd__o2bb2ai_1 _07190_ (.A1_N(_00810_),
    .A2_N(_00811_),
    .B1(_00840_),
    .B2(_00842_),
    .Y(_01033_));
 sky130_fd_sc_hd__o211ai_2 _07191_ (.A1(_00801_),
    .A2(_00809_),
    .B1(_00811_),
    .C1(_00843_),
    .Y(_01035_));
 sky130_fd_sc_hd__o2bb2ai_2 _07192_ (.A1_N(_00810_),
    .A2_N(_00811_),
    .B1(_00838_),
    .B2(_00839_),
    .Y(_01036_));
 sky130_fd_sc_hd__and4_2 _07193_ (.A(_00996_),
    .B(_01031_),
    .C(_01035_),
    .D(_01036_),
    .X(_01037_));
 sky130_fd_sc_hd__nand4_4 _07194_ (.A(_00996_),
    .B(_01031_),
    .C(_01035_),
    .D(_01036_),
    .Y(_01038_));
 sky130_fd_sc_hd__o2111ai_4 _07195_ (.A1(_01030_),
    .A2(_00995_),
    .B1(_00997_),
    .C1(_01032_),
    .D1(_01033_),
    .Y(_01039_));
 sky130_fd_sc_hd__o211ai_2 _07196_ (.A1(_00099_),
    .A2(_00451_),
    .B1(_00864_),
    .C1(_00865_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand4_2 _07197_ (.A(net32),
    .B(net2),
    .C(net37),
    .D(net36),
    .Y(_01041_));
 sky130_fd_sc_hd__nand2_1 _07198_ (.A(net31),
    .B(net38),
    .Y(_01042_));
 sky130_fd_sc_hd__a22oi_1 _07199_ (.A1(net32),
    .A2(net37),
    .B1(net36),
    .B2(net2),
    .Y(_01043_));
 sky130_fd_sc_hd__a22o_1 _07200_ (.A1(net32),
    .A2(net37),
    .B1(net36),
    .B2(net2),
    .X(_01044_));
 sky130_fd_sc_hd__and4_1 _07201_ (.A(_01044_),
    .B(net38),
    .C(net31),
    .D(_01041_),
    .X(_01046_));
 sky130_fd_sc_hd__o21ai_2 _07202_ (.A1(_01042_),
    .A2(_01043_),
    .B1(_01041_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand3_4 _07203_ (.A(_00866_),
    .B(_01040_),
    .C(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand2_1 _07204_ (.A(net29),
    .B(net39),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(net29),
    .B(net40),
    .Y(_01050_));
 sky130_fd_sc_hd__and4_2 _07206_ (.A(net30),
    .B(net29),
    .C(net39),
    .D(net40),
    .X(_01051_));
 sky130_fd_sc_hd__a22oi_2 _07207_ (.A1(net30),
    .A2(net39),
    .B1(net40),
    .B2(net29),
    .Y(_01052_));
 sky130_fd_sc_hd__a22o_1 _07208_ (.A1(net30),
    .A2(net39),
    .B1(net40),
    .B2(net29),
    .X(_01053_));
 sky130_fd_sc_hd__o2111a_2 _07209_ (.A1(_00861_),
    .A2(_01049_),
    .B1(net28),
    .C1(net41),
    .D1(_01053_),
    .X(_01054_));
 sky130_fd_sc_hd__o2111ai_4 _07210_ (.A1(_00861_),
    .A2(_01049_),
    .B1(net28),
    .C1(net41),
    .D1(_01053_),
    .Y(_01055_));
 sky130_fd_sc_hd__a31o_1 _07211_ (.A1(_01053_),
    .A2(net41),
    .A3(net28),
    .B1(_01051_),
    .X(_01057_));
 sky130_fd_sc_hd__a21o_2 _07212_ (.A1(_00866_),
    .A2(_01040_),
    .B1(_01047_),
    .X(_01058_));
 sky130_fd_sc_hd__o211a_1 _07213_ (.A1(_01051_),
    .A2(_01054_),
    .B1(_01058_),
    .C1(_01048_),
    .X(_01059_));
 sky130_fd_sc_hd__o211ai_4 _07214_ (.A1(_01051_),
    .A2(_01054_),
    .B1(_01058_),
    .C1(_01048_),
    .Y(_01060_));
 sky130_fd_sc_hd__a22oi_2 _07215_ (.A1(_00862_),
    .A2(_00866_),
    .B1(_00871_),
    .B2(_00860_),
    .Y(_01061_));
 sky130_fd_sc_hd__o21ai_1 _07216_ (.A1(_00859_),
    .A2(_00870_),
    .B1(_00868_),
    .Y(_01062_));
 sky130_fd_sc_hd__nor3_1 _07217_ (.A(_00868_),
    .B(_00870_),
    .C(_00859_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand3_1 _07218_ (.A(_00860_),
    .B(_00871_),
    .C(_00867_),
    .Y(_01064_));
 sky130_fd_sc_hd__o2bb2ai_4 _07219_ (.A1_N(_01048_),
    .A2_N(_01060_),
    .B1(_01061_),
    .B2(_01063_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand4_2 _07220_ (.A(_01048_),
    .B(_01060_),
    .C(_01062_),
    .D(_01064_),
    .Y(_01066_));
 sky130_fd_sc_hd__a22o_1 _07221_ (.A1(net26),
    .A2(net46),
    .B1(net47),
    .B2(net23),
    .X(_01068_));
 sky130_fd_sc_hd__nand4_2 _07222_ (.A(net26),
    .B(net23),
    .C(net46),
    .D(net47),
    .Y(_01069_));
 sky130_fd_sc_hd__a22o_1 _07223_ (.A1(_01068_),
    .A2(_01069_),
    .B1(net117),
    .B2(net12),
    .X(_01070_));
 sky130_fd_sc_hd__nand4_2 _07224_ (.A(net117),
    .B(_01068_),
    .C(_01069_),
    .D(net12),
    .Y(_01071_));
 sky130_fd_sc_hd__and2_1 _07225_ (.A(_01070_),
    .B(_01071_),
    .X(_01072_));
 sky130_fd_sc_hd__and4_1 _07226_ (.A(net28),
    .B(net27),
    .C(net43),
    .D(net42),
    .X(_01073_));
 sky130_fd_sc_hd__nand4_1 _07227_ (.A(net28),
    .B(net27),
    .C(net43),
    .D(net42),
    .Y(_01074_));
 sky130_fd_sc_hd__a22o_1 _07228_ (.A1(net27),
    .A2(net43),
    .B1(net42),
    .B2(net28),
    .X(_01075_));
 sky130_fd_sc_hd__and4_2 _07229_ (.A(_01075_),
    .B(net45),
    .C(net26),
    .D(_01074_),
    .X(_01076_));
 sky130_fd_sc_hd__a22o_1 _07230_ (.A1(net27),
    .A2(net45),
    .B1(_00887_),
    .B2(_00888_),
    .X(_01077_));
 sky130_fd_sc_hd__a211o_1 _07231_ (.A1(_00889_),
    .A2(_01077_),
    .B1(_01076_),
    .C1(_01073_),
    .X(_01079_));
 sky130_fd_sc_hd__o211a_1 _07232_ (.A1(_01073_),
    .A2(_01076_),
    .B1(_01077_),
    .C1(_00889_),
    .X(_01080_));
 sky130_fd_sc_hd__o211ai_2 _07233_ (.A1(_01073_),
    .A2(_01076_),
    .B1(_01077_),
    .C1(_00889_),
    .Y(_01081_));
 sky130_fd_sc_hd__and3_1 _07234_ (.A(_01072_),
    .B(_01079_),
    .C(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__nand4_2 _07235_ (.A(_01070_),
    .B(_01071_),
    .C(_01079_),
    .D(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _07236_ (.A1(_01079_),
    .A2(_01081_),
    .B1(_01072_),
    .Y(_01084_));
 sky130_fd_sc_hd__a22o_1 _07237_ (.A1(_01070_),
    .A2(_01071_),
    .B1(_01079_),
    .B2(_01081_),
    .X(_01085_));
 sky130_fd_sc_hd__nand4_4 _07238_ (.A(_01065_),
    .B(_01066_),
    .C(_01083_),
    .D(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _07239_ (.A(_01065_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__a21oi_2 _07240_ (.A1(_01018_),
    .A2(_01025_),
    .B1(_01022_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21o_1 _07241_ (.A1(_00878_),
    .A2(_00879_),
    .B1(_00899_),
    .X(_01090_));
 sky130_fd_sc_hd__nand3_1 _07242_ (.A(_00878_),
    .B(_00879_),
    .C(_00899_),
    .Y(_01091_));
 sky130_fd_sc_hd__a21o_1 _07243_ (.A1(_01090_),
    .A2(_01091_),
    .B1(_01088_),
    .X(_01092_));
 sky130_fd_sc_hd__nand3_1 _07244_ (.A(_01090_),
    .B(_01091_),
    .C(_01088_),
    .Y(_01093_));
 sky130_fd_sc_hd__a21oi_1 _07245_ (.A1(_01092_),
    .A2(_01093_),
    .B1(_01087_),
    .Y(_01094_));
 sky130_fd_sc_hd__a32o_1 _07246_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01088_),
    .B1(_01086_),
    .B2(_01065_),
    .X(_01095_));
 sky130_fd_sc_hd__and3_1 _07247_ (.A(_01087_),
    .B(_01092_),
    .C(_01093_),
    .X(_01096_));
 sky130_fd_sc_hd__and4_1 _07248_ (.A(_01065_),
    .B(_01086_),
    .C(_01092_),
    .D(_01093_),
    .X(_01097_));
 sky130_fd_sc_hd__a22oi_2 _07249_ (.A1(_01065_),
    .A2(_01086_),
    .B1(_01092_),
    .B2(_01093_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _07250_ (.A(_01094_),
    .B(_01096_),
    .Y(_01099_));
 sky130_fd_sc_hd__o21ai_2 _07251_ (.A1(_01097_),
    .A2(_01098_),
    .B1(_01039_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand3_2 _07252_ (.A(_00849_),
    .B(_00850_),
    .C(_00911_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _07253_ (.A(_00912_),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__a221oi_2 _07254_ (.A1(_01039_),
    .A2(_01099_),
    .B1(_01102_),
    .B2(_00912_),
    .C1(_01037_),
    .Y(_01104_));
 sky130_fd_sc_hd__a221o_1 _07255_ (.A1(_01039_),
    .A2(_01099_),
    .B1(_01102_),
    .B2(_00912_),
    .C1(_01037_),
    .X(_01105_));
 sky130_fd_sc_hd__a21oi_1 _07256_ (.A1(_01038_),
    .A2(_01101_),
    .B1(_01103_),
    .Y(_01106_));
 sky130_fd_sc_hd__a21o_1 _07257_ (.A1(_01038_),
    .A2(_01101_),
    .B1(_01103_),
    .X(_01107_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(_00883_),
    .B(_00885_),
    .Y(_01108_));
 sky130_fd_sc_hd__a2bb2oi_1 _07259_ (.A1_N(_00894_),
    .A2_N(_00896_),
    .B1(_01092_),
    .B2(_01095_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand4_1 _07260_ (.A(_00895_),
    .B(_00897_),
    .C(_01092_),
    .D(_01095_),
    .Y(_01110_));
 sky130_fd_sc_hd__and2b_1 _07261_ (.A_N(_01109_),
    .B(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _07262_ (.A(_01108_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__o21ai_2 _07263_ (.A1(_01104_),
    .A2(_01113_),
    .B1(_01107_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2b_1 _07264_ (.A_N(_00916_),
    .B(_00917_),
    .Y(_01115_));
 sky130_fd_sc_hd__xor2_1 _07265_ (.A(_00922_),
    .B(_01115_),
    .X(_01116_));
 sky130_fd_sc_hd__nor2_1 _07266_ (.A(_01114_),
    .B(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_01116_),
    .B(_01114_),
    .Y(_01118_));
 sky130_fd_sc_hd__a21o_1 _07268_ (.A1(_01112_),
    .A2(_01108_),
    .B1(_01109_),
    .X(_01119_));
 sky130_fd_sc_hd__inv_2 _07269_ (.A(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__a21oi_1 _07270_ (.A1(_01116_),
    .A2(_01114_),
    .B1(_01119_),
    .Y(_01121_));
 sky130_fd_sc_hd__o21ai_1 _07271_ (.A1(_01117_),
    .A2(_01120_),
    .B1(_01118_),
    .Y(_01123_));
 sky130_fd_sc_hd__xnor2_1 _07272_ (.A(_00939_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__and2b_1 _07273_ (.A_N(_01117_),
    .B(_01118_),
    .X(_01125_));
 sky130_fd_sc_hd__xor2_1 _07274_ (.A(_01120_),
    .B(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__nand2_2 _07275_ (.A(net11),
    .B(net33),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _07276_ (.A(net11),
    .B(net44),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(net10),
    .B(net55),
    .Y(_01129_));
 sky130_fd_sc_hd__a22oi_2 _07278_ (.A1(net11),
    .A2(net44),
    .B1(net33),
    .B2(net13),
    .Y(_01130_));
 sky130_fd_sc_hd__a22o_1 _07279_ (.A1(net11),
    .A2(net44),
    .B1(net33),
    .B2(net13),
    .X(_01131_));
 sky130_fd_sc_hd__nand3_1 _07280_ (.A(_01128_),
    .B(net33),
    .C(net13),
    .Y(_01132_));
 sky130_fd_sc_hd__nand3_1 _07281_ (.A(_00941_),
    .B(net44),
    .C(net11),
    .Y(_01134_));
 sky130_fd_sc_hd__o2111ai_4 _07282_ (.A1(_00942_),
    .A2(_01127_),
    .B1(net10),
    .C1(net55),
    .D1(_01131_),
    .Y(_01135_));
 sky130_fd_sc_hd__o22ai_4 _07283_ (.A1(_00942_),
    .A2(_01127_),
    .B1(_01129_),
    .B2(_01130_),
    .Y(_01136_));
 sky130_fd_sc_hd__o211ai_4 _07284_ (.A1(_00220_),
    .A2(_00341_),
    .B1(_00948_),
    .C1(_00949_),
    .Y(_01137_));
 sky130_fd_sc_hd__o31a_2 _07285_ (.A1(_00944_),
    .A2(_00945_),
    .A3(_00943_),
    .B1(_01136_),
    .X(_01138_));
 sky130_fd_sc_hd__nand3_2 _07286_ (.A(_00950_),
    .B(_01136_),
    .C(_01137_),
    .Y(_01139_));
 sky130_fd_sc_hd__a21oi_1 _07287_ (.A1(_00950_),
    .A2(_01137_),
    .B1(_01136_),
    .Y(_01140_));
 sky130_fd_sc_hd__a21o_2 _07288_ (.A1(_00950_),
    .A2(_01137_),
    .B1(_01136_),
    .X(_01141_));
 sky130_fd_sc_hd__nand2_1 _07289_ (.A(net8),
    .B(net60),
    .Y(_01142_));
 sky130_fd_sc_hd__a22oi_1 _07290_ (.A1(net10),
    .A2(net58),
    .B1(net59),
    .B2(net9),
    .Y(_01143_));
 sky130_fd_sc_hd__a22o_1 _07291_ (.A1(net10),
    .A2(net58),
    .B1(net59),
    .B2(net9),
    .X(_01145_));
 sky130_fd_sc_hd__nand4_2 _07292_ (.A(net9),
    .B(net10),
    .C(net58),
    .D(net59),
    .Y(_01146_));
 sky130_fd_sc_hd__and4_1 _07293_ (.A(_01145_),
    .B(_01146_),
    .C(net8),
    .D(net60),
    .X(_01147_));
 sky130_fd_sc_hd__o2bb2a_1 _07294_ (.A1_N(_01145_),
    .A2_N(_01146_),
    .B1(_00209_),
    .B2(_00352_),
    .X(_01148_));
 sky130_fd_sc_hd__a21o_1 _07295_ (.A1(_01145_),
    .A2(_01146_),
    .B1(_01142_),
    .X(_01149_));
 sky130_fd_sc_hd__o211ai_2 _07296_ (.A1(_00209_),
    .A2(_00352_),
    .B1(_01145_),
    .C1(_01146_),
    .Y(_01150_));
 sky130_fd_sc_hd__nand2_2 _07297_ (.A(_01149_),
    .B(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__a221oi_2 _07298_ (.A1(_01149_),
    .A2(_01150_),
    .B1(_01138_),
    .B2(_01137_),
    .C1(_01140_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand3_2 _07299_ (.A(_01139_),
    .B(_01141_),
    .C(_01151_),
    .Y(_01153_));
 sky130_fd_sc_hd__a22oi_4 _07300_ (.A1(_01137_),
    .A2(_01138_),
    .B1(_01141_),
    .B2(_01151_),
    .Y(_01154_));
 sky130_fd_sc_hd__a22o_1 _07301_ (.A1(_01137_),
    .A2(_01138_),
    .B1(_01141_),
    .B2(_01151_),
    .X(_01156_));
 sky130_fd_sc_hd__o211a_1 _07302_ (.A1(_00963_),
    .A2(_00965_),
    .B1(_00954_),
    .C1(_00955_),
    .X(_01157_));
 sky130_fd_sc_hd__o211ai_2 _07303_ (.A1(_00963_),
    .A2(_00965_),
    .B1(_00954_),
    .C1(_00955_),
    .Y(_01158_));
 sky130_fd_sc_hd__a21oi_2 _07304_ (.A1(_00954_),
    .A2(_00955_),
    .B1(_00967_),
    .Y(_01159_));
 sky130_fd_sc_hd__o2bb2ai_2 _07305_ (.A1_N(_00954_),
    .A2_N(_00955_),
    .B1(_00961_),
    .B2(_00962_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor3_2 _07306_ (.A(_01154_),
    .B(_01157_),
    .C(_01159_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand3_1 _07307_ (.A(_01156_),
    .B(_01158_),
    .C(_01160_),
    .Y(_01162_));
 sky130_fd_sc_hd__and4_1 _07308_ (.A(net7),
    .B(net6),
    .C(net62),
    .D(net61),
    .X(_01163_));
 sky130_fd_sc_hd__nand4_2 _07309_ (.A(net7),
    .B(net6),
    .C(net62),
    .D(net61),
    .Y(_01164_));
 sky130_fd_sc_hd__a22o_1 _07310_ (.A1(net6),
    .A2(net62),
    .B1(net61),
    .B2(net7),
    .X(_01165_));
 sky130_fd_sc_hd__and4_1 _07311_ (.A(_01165_),
    .B(net63),
    .C(net5),
    .D(_01164_),
    .X(_01167_));
 sky130_fd_sc_hd__nand4_2 _07312_ (.A(_01165_),
    .B(net63),
    .C(net5),
    .D(_01164_),
    .Y(_01168_));
 sky130_fd_sc_hd__o41a_1 _07313_ (.A1(_00176_),
    .A2(_00187_),
    .A3(_00374_),
    .A4(_00385_),
    .B1(_01168_),
    .X(_01169_));
 sky130_fd_sc_hd__o21ai_2 _07314_ (.A1(_01142_),
    .A2(_01143_),
    .B1(_01146_),
    .Y(_01170_));
 sky130_fd_sc_hd__o2bb2ai_1 _07315_ (.A1_N(_00974_),
    .A2_N(_00975_),
    .B1(_00187_),
    .B2(_00396_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand3_2 _07316_ (.A(_00976_),
    .B(_01170_),
    .C(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__a21oi_1 _07317_ (.A1(_00976_),
    .A2(_01171_),
    .B1(_01170_),
    .Y(_01173_));
 sky130_fd_sc_hd__a21o_1 _07318_ (.A1(_00976_),
    .A2(_01171_),
    .B1(_01170_),
    .X(_01174_));
 sky130_fd_sc_hd__o211a_1 _07319_ (.A1(_01163_),
    .A2(_01167_),
    .B1(_01172_),
    .C1(_01174_),
    .X(_01175_));
 sky130_fd_sc_hd__a21boi_2 _07320_ (.A1(_01172_),
    .A2(_01174_),
    .B1_N(_01169_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _07321_ (.A(_01175_),
    .B(_01176_),
    .Y(_01178_));
 sky130_fd_sc_hd__a21oi_4 _07322_ (.A1(_01158_),
    .A2(_01160_),
    .B1(_01156_),
    .Y(_01179_));
 sky130_fd_sc_hd__o21ai_1 _07323_ (.A1(_01157_),
    .A2(_01159_),
    .B1(_01154_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(_01178_),
    .B(_01162_),
    .Y(_01181_));
 sky130_fd_sc_hd__and3_1 _07325_ (.A(_01178_),
    .B(_01180_),
    .C(_01162_),
    .X(_01182_));
 sky130_fd_sc_hd__nand3_1 _07326_ (.A(_01178_),
    .B(_01180_),
    .C(_01162_),
    .Y(_01183_));
 sky130_fd_sc_hd__o32a_2 _07327_ (.A1(_01154_),
    .A2(_01157_),
    .A3(_01159_),
    .B1(_01179_),
    .B2(_01181_),
    .X(_01184_));
 sky130_fd_sc_hd__o211ai_4 _07328_ (.A1(_00985_),
    .A2(_00986_),
    .B1(_00972_),
    .C1(_00973_),
    .Y(_01185_));
 sky130_fd_sc_hd__o2bb2ai_2 _07329_ (.A1_N(_00972_),
    .A2_N(_00973_),
    .B1(_00987_),
    .B2(_00988_),
    .Y(_01186_));
 sky130_fd_sc_hd__o211ai_2 _07330_ (.A1(_00987_),
    .A2(_00988_),
    .B1(_00972_),
    .C1(_00973_),
    .Y(_01187_));
 sky130_fd_sc_hd__o2bb2ai_2 _07331_ (.A1_N(_00972_),
    .A2_N(_00973_),
    .B1(_00985_),
    .B2(_00986_),
    .Y(_01189_));
 sky130_fd_sc_hd__o211a_2 _07332_ (.A1(_01161_),
    .A2(_01182_),
    .B1(_01187_),
    .C1(_01189_),
    .X(_01190_));
 sky130_fd_sc_hd__o211ai_4 _07333_ (.A1(_01161_),
    .A2(_01182_),
    .B1(_01187_),
    .C1(_01189_),
    .Y(_01191_));
 sky130_fd_sc_hd__and4_1 _07334_ (.A(net3),
    .B(net4),
    .C(net64),
    .D(net34),
    .X(_01192_));
 sky130_fd_sc_hd__nand4_1 _07335_ (.A(net3),
    .B(net4),
    .C(net64),
    .D(net34),
    .Y(_01193_));
 sky130_fd_sc_hd__a22oi_4 _07336_ (.A1(net4),
    .A2(net64),
    .B1(net34),
    .B2(net3),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _07337_ (.A(net2),
    .B(net35),
    .Y(_01195_));
 sky130_fd_sc_hd__nand4b_2 _07338_ (.A_N(_01194_),
    .B(net35),
    .C(net2),
    .D(_01193_),
    .Y(_01196_));
 sky130_fd_sc_hd__o21ai_1 _07339_ (.A1(_01195_),
    .A2(_01194_),
    .B1(_01193_),
    .Y(_01197_));
 sky130_fd_sc_hd__o211ai_2 _07340_ (.A1(_00132_),
    .A2(_00407_),
    .B1(_01003_),
    .C1(_01004_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand3_1 _07341_ (.A(_01005_),
    .B(_01197_),
    .C(_01198_),
    .Y(_01200_));
 sky130_fd_sc_hd__a21oi_1 _07342_ (.A1(_01005_),
    .A2(_01198_),
    .B1(_01197_),
    .Y(_01201_));
 sky130_fd_sc_hd__a21o_1 _07343_ (.A1(_01005_),
    .A2(_01198_),
    .B1(_01197_),
    .X(_01202_));
 sky130_fd_sc_hd__a22oi_2 _07344_ (.A1(net31),
    .A2(net38),
    .B1(_01041_),
    .B2(_01044_),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_1 _07345_ (.A(_01046_),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__o31a_2 _07346_ (.A1(_01046_),
    .A2(_01201_),
    .A3(_01203_),
    .B1(_01200_),
    .X(_01205_));
 sky130_fd_sc_hd__o21ai_2 _07347_ (.A1(_01169_),
    .A2(_01173_),
    .B1(_01172_),
    .Y(_01206_));
 sky130_fd_sc_hd__o22ai_2 _07348_ (.A1(_00856_),
    .A2(_01011_),
    .B1(_01014_),
    .B2(_01010_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand3_1 _07349_ (.A(_01016_),
    .B(_01206_),
    .C(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__a21oi_1 _07350_ (.A1(_01016_),
    .A2(_01207_),
    .B1(_01206_),
    .Y(_01209_));
 sky130_fd_sc_hd__a21o_1 _07351_ (.A1(_01016_),
    .A2(_01207_),
    .B1(_01206_),
    .X(_01211_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(_01208_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__xor2_1 _07353_ (.A(_01205_),
    .B(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__xnor2_2 _07354_ (.A(_01205_),
    .B(_01212_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand3_2 _07355_ (.A(_01186_),
    .B(_01184_),
    .C(_01185_),
    .Y(_01215_));
 sky130_fd_sc_hd__a31oi_4 _07356_ (.A1(_01186_),
    .A2(_01184_),
    .A3(_01185_),
    .B1(_01214_),
    .Y(_01216_));
 sky130_fd_sc_hd__a31o_2 _07357_ (.A1(_01186_),
    .A2(_01184_),
    .A3(_01185_),
    .B1(_01214_),
    .X(_01217_));
 sky130_fd_sc_hd__a21oi_1 _07358_ (.A1(_01213_),
    .A2(_01215_),
    .B1(_01190_),
    .Y(_01218_));
 sky130_fd_sc_hd__o211ai_4 _07359_ (.A1(_01026_),
    .A2(_01027_),
    .B1(_00996_),
    .C1(_00997_),
    .Y(_01219_));
 sky130_fd_sc_hd__o2bb2ai_2 _07360_ (.A1_N(_00996_),
    .A2_N(_00997_),
    .B1(_01028_),
    .B2(_01029_),
    .Y(_01220_));
 sky130_fd_sc_hd__o211ai_2 _07361_ (.A1(_01028_),
    .A2(_01029_),
    .B1(_00996_),
    .C1(_00997_),
    .Y(_01222_));
 sky130_fd_sc_hd__o2bb2ai_2 _07362_ (.A1_N(_00996_),
    .A2_N(_00997_),
    .B1(_01026_),
    .B2(_01027_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand4_4 _07363_ (.A(_01191_),
    .B(_01217_),
    .C(_01219_),
    .D(_01220_),
    .Y(_01224_));
 sky130_fd_sc_hd__o211a_1 _07364_ (.A1(_01190_),
    .A2(_01216_),
    .B1(_01222_),
    .C1(_01223_),
    .X(_01225_));
 sky130_fd_sc_hd__o211ai_4 _07365_ (.A1(_01190_),
    .A2(_01216_),
    .B1(_01222_),
    .C1(_01223_),
    .Y(_01226_));
 sky130_fd_sc_hd__and4_1 _07366_ (.A(net32),
    .B(net31),
    .C(net37),
    .D(net36),
    .X(_01227_));
 sky130_fd_sc_hd__nand4_1 _07367_ (.A(net32),
    .B(net31),
    .C(net37),
    .D(net36),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(net30),
    .B(net38),
    .Y(_01229_));
 sky130_fd_sc_hd__a22oi_2 _07369_ (.A1(net31),
    .A2(net37),
    .B1(net36),
    .B2(net32),
    .Y(_01230_));
 sky130_fd_sc_hd__a22o_1 _07370_ (.A1(net31),
    .A2(net37),
    .B1(net36),
    .B2(net32),
    .X(_01231_));
 sky130_fd_sc_hd__and4_2 _07371_ (.A(_01231_),
    .B(net38),
    .C(net30),
    .D(_01228_),
    .X(_01233_));
 sky130_fd_sc_hd__or3_2 _07372_ (.A(_01229_),
    .B(_01230_),
    .C(_01227_),
    .X(_01234_));
 sky130_fd_sc_hd__o21ai_1 _07373_ (.A1(_01229_),
    .A2(_01230_),
    .B1(_01228_),
    .Y(_01235_));
 sky130_fd_sc_hd__o22a_1 _07374_ (.A1(_00066_),
    .A2(_00451_),
    .B1(_01051_),
    .B2(_01052_),
    .X(_01236_));
 sky130_fd_sc_hd__o22ai_2 _07375_ (.A1(_00066_),
    .A2(_00451_),
    .B1(_01051_),
    .B2(_01052_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_01055_),
    .B(_01235_),
    .Y(_01238_));
 sky130_fd_sc_hd__and3_2 _07377_ (.A(_01055_),
    .B(_01235_),
    .C(_01237_),
    .X(_01239_));
 sky130_fd_sc_hd__o211ai_4 _07378_ (.A1(_01227_),
    .A2(_01233_),
    .B1(_01237_),
    .C1(_01055_),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _07379_ (.A(net28),
    .B(net39),
    .Y(_01241_));
 sky130_fd_sc_hd__and4_2 _07380_ (.A(net28),
    .B(net29),
    .C(net39),
    .D(net40),
    .X(_01242_));
 sky130_fd_sc_hd__nand4_1 _07381_ (.A(net28),
    .B(net29),
    .C(net39),
    .D(net40),
    .Y(_01244_));
 sky130_fd_sc_hd__a22o_1 _07382_ (.A1(net29),
    .A2(net39),
    .B1(net40),
    .B2(net28),
    .X(_01245_));
 sky130_fd_sc_hd__and2_1 _07383_ (.A(net27),
    .B(net41),
    .X(_01246_));
 sky130_fd_sc_hd__o211a_2 _07384_ (.A1(_01050_),
    .A2(_01241_),
    .B1(_01246_),
    .C1(_01245_),
    .X(_01247_));
 sky130_fd_sc_hd__o2111ai_2 _07385_ (.A1(_01050_),
    .A2(_01241_),
    .B1(net27),
    .C1(net41),
    .D1(_01245_),
    .Y(_01248_));
 sky130_fd_sc_hd__a31o_1 _07386_ (.A1(_01245_),
    .A2(net41),
    .A3(net27),
    .B1(_01242_),
    .X(_01249_));
 sky130_fd_sc_hd__o21bai_4 _07387_ (.A1(_01054_),
    .A2(_01236_),
    .B1_N(_01235_),
    .Y(_01250_));
 sky130_fd_sc_hd__o21a_1 _07388_ (.A1(_01242_),
    .A2(_01247_),
    .B1(_01250_),
    .X(_01251_));
 sky130_fd_sc_hd__o21ai_4 _07389_ (.A1(_01242_),
    .A2(_01247_),
    .B1(_01250_),
    .Y(_01252_));
 sky130_fd_sc_hd__o221a_1 _07390_ (.A1(_01236_),
    .A2(_01238_),
    .B1(_01242_),
    .B2(_01247_),
    .C1(_01250_),
    .X(_01253_));
 sky130_fd_sc_hd__a21oi_1 _07391_ (.A1(_01048_),
    .A2(_01058_),
    .B1(_01057_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21o_1 _07392_ (.A1(_01048_),
    .A2(_01058_),
    .B1(_01057_),
    .X(_01256_));
 sky130_fd_sc_hd__o211ai_4 _07393_ (.A1(_01239_),
    .A2(_01251_),
    .B1(_01256_),
    .C1(_01060_),
    .Y(_01257_));
 sky130_fd_sc_hd__a22o_1 _07394_ (.A1(net23),
    .A2(net46),
    .B1(net47),
    .B2(net12),
    .X(_01258_));
 sky130_fd_sc_hd__nand4_4 _07395_ (.A(net12),
    .B(net23),
    .C(net46),
    .D(net47),
    .Y(_01259_));
 sky130_fd_sc_hd__a22o_1 _07396_ (.A1(_01258_),
    .A2(_01259_),
    .B1(net117),
    .B2(net1),
    .X(_01260_));
 sky130_fd_sc_hd__nand4_4 _07397_ (.A(net117),
    .B(_01258_),
    .C(_01259_),
    .D(net1),
    .Y(_01261_));
 sky130_fd_sc_hd__nand4_4 _07398_ (.A(net26),
    .B(net27),
    .C(net43),
    .D(net42),
    .Y(_01262_));
 sky130_fd_sc_hd__a22o_1 _07399_ (.A1(net26),
    .A2(net43),
    .B1(net42),
    .B2(net27),
    .X(_01263_));
 sky130_fd_sc_hd__nand4_4 _07400_ (.A(_01263_),
    .B(net45),
    .C(net23),
    .D(_01262_),
    .Y(_01264_));
 sky130_fd_sc_hd__a22oi_2 _07401_ (.A1(net26),
    .A2(net45),
    .B1(_01074_),
    .B2(_01075_),
    .Y(_01266_));
 sky130_fd_sc_hd__o211ai_2 _07402_ (.A1(_01076_),
    .A2(_01266_),
    .B1(_01264_),
    .C1(_01262_),
    .Y(_01267_));
 sky130_fd_sc_hd__a211o_2 _07403_ (.A1(_01262_),
    .A2(_01264_),
    .B1(_01266_),
    .C1(_01076_),
    .X(_01268_));
 sky130_fd_sc_hd__nand4_4 _07404_ (.A(_01260_),
    .B(_01261_),
    .C(_01267_),
    .D(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__a22o_1 _07405_ (.A1(_01260_),
    .A2(_01261_),
    .B1(_01267_),
    .B2(_01268_),
    .X(_01270_));
 sky130_fd_sc_hd__o211ai_4 _07406_ (.A1(_01059_),
    .A2(_01255_),
    .B1(_01252_),
    .C1(_01240_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand4_4 _07407_ (.A(_01257_),
    .B(_01269_),
    .C(_01270_),
    .D(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_01257_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__o21ai_2 _07409_ (.A1(_01205_),
    .A2(_01209_),
    .B1(_01208_),
    .Y(_01274_));
 sky130_fd_sc_hd__o2bb2ai_1 _07410_ (.A1_N(_01065_),
    .A2_N(_01066_),
    .B1(_01082_),
    .B2(_01084_),
    .Y(_01275_));
 sky130_fd_sc_hd__a21oi_2 _07411_ (.A1(_01086_),
    .A2(_01275_),
    .B1(_01274_),
    .Y(_01277_));
 sky130_fd_sc_hd__a21o_1 _07412_ (.A1(_01086_),
    .A2(_01275_),
    .B1(_01274_),
    .X(_01278_));
 sky130_fd_sc_hd__and3_2 _07413_ (.A(_01086_),
    .B(_01274_),
    .C(_01275_),
    .X(_01279_));
 sky130_fd_sc_hd__a211oi_2 _07414_ (.A1(_01257_),
    .A2(_01272_),
    .B1(_01277_),
    .C1(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__a211o_1 _07415_ (.A1(_01257_),
    .A2(_01272_),
    .B1(_01277_),
    .C1(_01279_),
    .X(_01281_));
 sky130_fd_sc_hd__o211a_1 _07416_ (.A1(_01277_),
    .A2(_01279_),
    .B1(_01257_),
    .C1(_01272_),
    .X(_01282_));
 sky130_fd_sc_hd__o211ai_2 _07417_ (.A1(_01277_),
    .A2(_01279_),
    .B1(_01257_),
    .C1(_01272_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_2 _07418_ (.A(_01281_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__a31oi_2 _07419_ (.A1(_01218_),
    .A2(_01219_),
    .A3(_01220_),
    .B1(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__a31o_1 _07420_ (.A1(_01218_),
    .A2(_01219_),
    .A3(_01220_),
    .B1(_01284_),
    .X(_01286_));
 sky130_fd_sc_hd__a21o_1 _07421_ (.A1(_01038_),
    .A2(_01039_),
    .B1(_01099_),
    .X(_01288_));
 sky130_fd_sc_hd__o2bb2ai_1 _07422_ (.A1_N(_01038_),
    .A2_N(_01039_),
    .B1(_01097_),
    .B2(_01098_),
    .Y(_01289_));
 sky130_fd_sc_hd__o211ai_1 _07423_ (.A1(_01094_),
    .A2(_01096_),
    .B1(_01038_),
    .C1(_01039_),
    .Y(_01290_));
 sky130_fd_sc_hd__o221ai_4 _07424_ (.A1(_01037_),
    .A2(_01101_),
    .B1(_01225_),
    .B2(_01285_),
    .C1(_01288_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand4_2 _07425_ (.A(_01226_),
    .B(_01286_),
    .C(_01289_),
    .D(_01290_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(_01069_),
    .B(_01071_),
    .Y(_01293_));
 sky130_fd_sc_hd__a31o_1 _07427_ (.A1(_01070_),
    .A2(_01071_),
    .A3(_01079_),
    .B1(_01080_),
    .X(_01294_));
 sky130_fd_sc_hd__o22ai_1 _07428_ (.A1(_01080_),
    .A2(_01082_),
    .B1(_01279_),
    .B2(_01280_),
    .Y(_01295_));
 sky130_fd_sc_hd__a211o_1 _07429_ (.A1(_01273_),
    .A2(_01278_),
    .B1(_01279_),
    .C1(_01294_),
    .X(_01296_));
 sky130_fd_sc_hd__nand2_1 _07430_ (.A(_01295_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(_01293_),
    .B(_01297_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _07432_ (.A(_01299_),
    .B(_01292_),
    .Y(_01300_));
 sky130_fd_sc_hd__o21bai_1 _07433_ (.A1(_01104_),
    .A2(_01106_),
    .B1_N(_01113_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand3_1 _07434_ (.A(_01105_),
    .B(_01107_),
    .C(_01113_),
    .Y(_01302_));
 sky130_fd_sc_hd__and4_1 _07435_ (.A(_01291_),
    .B(_01300_),
    .C(_01301_),
    .D(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__a22oi_2 _07436_ (.A1(_01291_),
    .A2(_01300_),
    .B1(_01301_),
    .B2(_01302_),
    .Y(_01304_));
 sky130_fd_sc_hd__a21boi_1 _07437_ (.A1(_01293_),
    .A2(_01296_),
    .B1_N(_01295_),
    .Y(_01305_));
 sky130_fd_sc_hd__o21ba_1 _07438_ (.A1(_01303_),
    .A2(_01305_),
    .B1_N(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__nor3_1 _07439_ (.A(_01303_),
    .B(_01304_),
    .C(_01305_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _07440_ (.A(_01126_),
    .B(_01306_),
    .Y(_01308_));
 sky130_fd_sc_hd__or2_1 _07441_ (.A(_01306_),
    .B(_01126_),
    .X(_01310_));
 sky130_fd_sc_hd__o21a_1 _07442_ (.A1(_01303_),
    .A2(_01304_),
    .B1(_01305_),
    .X(_01311_));
 sky130_fd_sc_hd__nor2_2 _07443_ (.A(_01307_),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__o22ai_4 _07444_ (.A1(_01175_),
    .A2(_01176_),
    .B1(_01179_),
    .B2(_01161_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _07445_ (.A(net10),
    .B(net33),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(net10),
    .B(net44),
    .Y(_01315_));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(net9),
    .B(net55),
    .Y(_01316_));
 sky130_fd_sc_hd__a22oi_1 _07448_ (.A1(net10),
    .A2(net44),
    .B1(net33),
    .B2(net11),
    .Y(_01317_));
 sky130_fd_sc_hd__a22o_1 _07449_ (.A1(net10),
    .A2(net44),
    .B1(net33),
    .B2(net11),
    .X(_01318_));
 sky130_fd_sc_hd__nand3_1 _07450_ (.A(_01315_),
    .B(net33),
    .C(net11),
    .Y(_01319_));
 sky130_fd_sc_hd__nand3_1 _07451_ (.A(_01127_),
    .B(net44),
    .C(net10),
    .Y(_01321_));
 sky130_fd_sc_hd__o2111ai_2 _07452_ (.A1(_01128_),
    .A2(_01314_),
    .B1(net9),
    .C1(net55),
    .D1(_01318_),
    .Y(_01322_));
 sky130_fd_sc_hd__o22ai_2 _07453_ (.A1(_01128_),
    .A2(_01314_),
    .B1(_01316_),
    .B2(_01317_),
    .Y(_01323_));
 sky130_fd_sc_hd__and3_1 _07454_ (.A(_01129_),
    .B(_01132_),
    .C(_01134_),
    .X(_01324_));
 sky130_fd_sc_hd__o211ai_2 _07455_ (.A1(_00231_),
    .A2(_00341_),
    .B1(_01132_),
    .C1(_01134_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _07456_ (.A(_01135_),
    .B(_01323_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand3_2 _07457_ (.A(_01135_),
    .B(_01323_),
    .C(_01325_),
    .Y(_01327_));
 sky130_fd_sc_hd__a21o_2 _07458_ (.A1(_01135_),
    .A2(_01325_),
    .B1(_01323_),
    .X(_01328_));
 sky130_fd_sc_hd__nand2_1 _07459_ (.A(net7),
    .B(net60),
    .Y(_01329_));
 sky130_fd_sc_hd__a22oi_1 _07460_ (.A1(net9),
    .A2(net58),
    .B1(net59),
    .B2(net8),
    .Y(_01330_));
 sky130_fd_sc_hd__a22o_1 _07461_ (.A1(net9),
    .A2(net58),
    .B1(net59),
    .B2(net8),
    .X(_01332_));
 sky130_fd_sc_hd__and4_1 _07462_ (.A(net9),
    .B(net8),
    .C(net58),
    .D(net59),
    .X(_01333_));
 sky130_fd_sc_hd__nand4_2 _07463_ (.A(net9),
    .B(net8),
    .C(net58),
    .D(net59),
    .Y(_01334_));
 sky130_fd_sc_hd__and4_1 _07464_ (.A(_01332_),
    .B(_01334_),
    .C(net7),
    .D(net60),
    .X(_01335_));
 sky130_fd_sc_hd__o22a_1 _07465_ (.A1(_00176_),
    .A2(_00352_),
    .B1(_01330_),
    .B2(_01333_),
    .X(_01336_));
 sky130_fd_sc_hd__o211a_1 _07466_ (.A1(_01330_),
    .A2(_01333_),
    .B1(net7),
    .C1(net60),
    .X(_01337_));
 sky130_fd_sc_hd__a21o_1 _07467_ (.A1(_01332_),
    .A2(_01334_),
    .B1(_01329_),
    .X(_01338_));
 sky130_fd_sc_hd__and3_1 _07468_ (.A(_01329_),
    .B(_01332_),
    .C(_01334_),
    .X(_01339_));
 sky130_fd_sc_hd__o211ai_1 _07469_ (.A1(_00176_),
    .A2(_00352_),
    .B1(_01332_),
    .C1(_01334_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(_01338_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o221a_2 _07471_ (.A1(_01324_),
    .A2(_01326_),
    .B1(_01337_),
    .B2(_01339_),
    .C1(_01328_),
    .X(_01343_));
 sky130_fd_sc_hd__o221ai_4 _07472_ (.A1(_01324_),
    .A2(_01326_),
    .B1(_01337_),
    .B2(_01339_),
    .C1(_01328_),
    .Y(_01344_));
 sky130_fd_sc_hd__a21boi_1 _07473_ (.A1(_01328_),
    .A2(_01341_),
    .B1_N(_01327_),
    .Y(_01345_));
 sky130_fd_sc_hd__a2bb2o_1 _07474_ (.A1_N(_01324_),
    .A2_N(_01326_),
    .B1(_01341_),
    .B2(_01328_),
    .X(_01346_));
 sky130_fd_sc_hd__a21oi_1 _07475_ (.A1(_01139_),
    .A2(_01141_),
    .B1(_01151_),
    .Y(_01347_));
 sky130_fd_sc_hd__o2bb2ai_2 _07476_ (.A1_N(_01139_),
    .A2_N(_01141_),
    .B1(_01147_),
    .B2(_01148_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21oi_4 _07477_ (.A1(_01153_),
    .A2(_01348_),
    .B1(_01346_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor3_1 _07478_ (.A(_01152_),
    .B(_01345_),
    .C(_01347_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand3_2 _07479_ (.A(_01153_),
    .B(_01346_),
    .C(_01348_),
    .Y(_01351_));
 sky130_fd_sc_hd__a31o_1 _07480_ (.A1(_01332_),
    .A2(net60),
    .A3(net7),
    .B1(_01333_),
    .X(_01352_));
 sky130_fd_sc_hd__o2bb2ai_1 _07481_ (.A1_N(_01164_),
    .A2_N(_01165_),
    .B1(_00154_),
    .B2(_00396_),
    .Y(_01354_));
 sky130_fd_sc_hd__a21oi_1 _07482_ (.A1(_01168_),
    .A2(_01354_),
    .B1(_01352_),
    .Y(_01355_));
 sky130_fd_sc_hd__a21o_1 _07483_ (.A1(_01168_),
    .A2(_01354_),
    .B1(_01352_),
    .X(_01356_));
 sky130_fd_sc_hd__o211ai_2 _07484_ (.A1(_01333_),
    .A2(_01335_),
    .B1(_01354_),
    .C1(_01168_),
    .Y(_01357_));
 sky130_fd_sc_hd__a22oi_1 _07485_ (.A1(net5),
    .A2(net62),
    .B1(net61),
    .B2(net6),
    .Y(_01358_));
 sky130_fd_sc_hd__a22o_1 _07486_ (.A1(net5),
    .A2(net62),
    .B1(net61),
    .B2(net6),
    .X(_01359_));
 sky130_fd_sc_hd__nand2_1 _07487_ (.A(net5),
    .B(net61),
    .Y(_01360_));
 sky130_fd_sc_hd__nand4_4 _07488_ (.A(net5),
    .B(net6),
    .C(net62),
    .D(net61),
    .Y(_01361_));
 sky130_fd_sc_hd__o32a_1 _07489_ (.A1(_00187_),
    .A2(_00374_),
    .A3(_01360_),
    .B1(_00396_),
    .B2(_00165_),
    .X(_01362_));
 sky130_fd_sc_hd__o31a_1 _07490_ (.A1(_00165_),
    .A2(_00396_),
    .A3(_01358_),
    .B1(_01361_),
    .X(_01363_));
 sky130_fd_sc_hd__nand3b_1 _07491_ (.A_N(_01363_),
    .B(_01357_),
    .C(_01356_),
    .Y(_01365_));
 sky130_fd_sc_hd__o2bb2ai_1 _07492_ (.A1_N(_01356_),
    .A2_N(_01357_),
    .B1(_01358_),
    .B2(_01362_),
    .Y(_01366_));
 sky130_fd_sc_hd__nand2_2 _07493_ (.A(_01365_),
    .B(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__o31a_1 _07494_ (.A1(_01152_),
    .A2(_01345_),
    .A3(_01347_),
    .B1(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__o21ai_2 _07495_ (.A1(_01367_),
    .A2(_01349_),
    .B1(_01351_),
    .Y(_01369_));
 sky130_fd_sc_hd__o211a_1 _07496_ (.A1(_01179_),
    .A2(_01181_),
    .B1(_01313_),
    .C1(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__o211ai_4 _07497_ (.A1(_01179_),
    .A2(_01181_),
    .B1(_01313_),
    .C1(_01369_),
    .Y(_01371_));
 sky130_fd_sc_hd__o21ai_1 _07498_ (.A1(_01363_),
    .A2(_01355_),
    .B1(_01357_),
    .Y(_01372_));
 sky130_fd_sc_hd__o2bb2ai_1 _07499_ (.A1_N(_01200_),
    .A2_N(_01202_),
    .B1(_01203_),
    .B2(_01046_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand3_1 _07500_ (.A(_01204_),
    .B(_01202_),
    .C(_01200_),
    .Y(_01374_));
 sky130_fd_sc_hd__a21o_1 _07501_ (.A1(_01373_),
    .A2(_01374_),
    .B1(_01372_),
    .X(_01376_));
 sky130_fd_sc_hd__nand3_1 _07502_ (.A(_01372_),
    .B(_01373_),
    .C(_01374_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _07503_ (.A(net2),
    .B(net64),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_2 _07504_ (.A(net2),
    .B(net34),
    .Y(_01379_));
 sky130_fd_sc_hd__and4_1 _07505_ (.A(net3),
    .B(net2),
    .C(net64),
    .D(net34),
    .X(_01380_));
 sky130_fd_sc_hd__a22o_1 _07506_ (.A1(net3),
    .A2(net64),
    .B1(net34),
    .B2(net2),
    .X(_01381_));
 sky130_fd_sc_hd__nand3_1 _07507_ (.A(_01379_),
    .B(net64),
    .C(net3),
    .Y(_01382_));
 sky130_fd_sc_hd__a21o_1 _07508_ (.A1(net3),
    .A2(net64),
    .B1(_01379_),
    .X(_01383_));
 sky130_fd_sc_hd__nand4b_2 _07509_ (.A_N(_01380_),
    .B(_01381_),
    .C(net32),
    .D(net35),
    .Y(_01384_));
 sky130_fd_sc_hd__a31o_1 _07510_ (.A1(_01381_),
    .A2(net35),
    .A3(net32),
    .B1(_01380_),
    .X(_01385_));
 sky130_fd_sc_hd__o22ai_4 _07511_ (.A1(_00143_),
    .A2(_00407_),
    .B1(_01192_),
    .B2(_01194_),
    .Y(_01387_));
 sky130_fd_sc_hd__and3_1 _07512_ (.A(_01196_),
    .B(_01385_),
    .C(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__nand3_2 _07513_ (.A(_01196_),
    .B(_01385_),
    .C(_01387_),
    .Y(_01389_));
 sky130_fd_sc_hd__a21o_1 _07514_ (.A1(_01196_),
    .A2(_01387_),
    .B1(_01385_),
    .X(_01390_));
 sky130_fd_sc_hd__o2bb2a_1 _07515_ (.A1_N(net30),
    .A2_N(net38),
    .B1(_01227_),
    .B2(_01230_),
    .X(_01391_));
 sky130_fd_sc_hd__a22o_1 _07516_ (.A1(net30),
    .A2(net38),
    .B1(_01228_),
    .B2(_01231_),
    .X(_01392_));
 sky130_fd_sc_hd__a31o_1 _07517_ (.A1(_01234_),
    .A2(_01390_),
    .A3(_01392_),
    .B1(_01388_),
    .X(_01393_));
 sky130_fd_sc_hd__and3_1 _07518_ (.A(_01376_),
    .B(_01377_),
    .C(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__a21oi_2 _07519_ (.A1(_01376_),
    .A2(_01377_),
    .B1(_01393_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_1 _07520_ (.A(_01394_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__a21oi_2 _07521_ (.A1(_01183_),
    .A2(_01313_),
    .B1(_01369_),
    .Y(_01398_));
 sky130_fd_sc_hd__o2bb2ai_2 _07522_ (.A1_N(_01183_),
    .A2_N(_01313_),
    .B1(_01349_),
    .B2(_01368_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand3_4 _07523_ (.A(_01396_),
    .B(_01399_),
    .C(_01371_),
    .Y(_01400_));
 sky130_fd_sc_hd__o31a_1 _07524_ (.A1(_01394_),
    .A2(_01395_),
    .A3(_01398_),
    .B1(_01371_),
    .X(_01401_));
 sky130_fd_sc_hd__a21o_1 _07525_ (.A1(_01396_),
    .A2(_01399_),
    .B1(_01370_),
    .X(_01402_));
 sky130_fd_sc_hd__a21oi_1 _07526_ (.A1(_01191_),
    .A2(_01215_),
    .B1(_01213_),
    .Y(_01403_));
 sky130_fd_sc_hd__a21o_1 _07527_ (.A1(_01191_),
    .A2(_01215_),
    .B1(_01213_),
    .X(_01404_));
 sky130_fd_sc_hd__nand3_1 _07528_ (.A(_01191_),
    .B(_01214_),
    .C(_01215_),
    .Y(_01405_));
 sky130_fd_sc_hd__a21o_1 _07529_ (.A1(_01191_),
    .A2(_01215_),
    .B1(_01214_),
    .X(_01406_));
 sky130_fd_sc_hd__nand3_4 _07530_ (.A(_01406_),
    .B(_01401_),
    .C(_01405_),
    .Y(_01407_));
 sky130_fd_sc_hd__a221oi_4 _07531_ (.A1(_01191_),
    .A2(_01216_),
    .B1(_01371_),
    .B2(_01400_),
    .C1(_01403_),
    .Y(_01409_));
 sky130_fd_sc_hd__o211ai_4 _07532_ (.A1(_01190_),
    .A2(_01217_),
    .B1(_01402_),
    .C1(_01404_),
    .Y(_01410_));
 sky130_fd_sc_hd__a21bo_1 _07533_ (.A1(_01376_),
    .A2(_01393_),
    .B1_N(_01377_),
    .X(_01411_));
 sky130_fd_sc_hd__a22o_1 _07534_ (.A1(_01269_),
    .A2(_01270_),
    .B1(_01271_),
    .B2(_01257_),
    .X(_01412_));
 sky130_fd_sc_hd__a21oi_1 _07535_ (.A1(_01272_),
    .A2(_01412_),
    .B1(_01411_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21o_1 _07536_ (.A1(_01272_),
    .A2(_01412_),
    .B1(_01411_),
    .X(_01414_));
 sky130_fd_sc_hd__nand3_2 _07537_ (.A(_01272_),
    .B(_01411_),
    .C(_01412_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21oi_1 _07538_ (.A1(_01240_),
    .A2(_01250_),
    .B1(_01249_),
    .Y(_01416_));
 sky130_fd_sc_hd__a21o_1 _07539_ (.A1(_01240_),
    .A2(_01250_),
    .B1(_01249_),
    .X(_01417_));
 sky130_fd_sc_hd__and4_1 _07540_ (.A(net30),
    .B(net31),
    .C(net37),
    .D(net36),
    .X(_01418_));
 sky130_fd_sc_hd__nand4_1 _07541_ (.A(net30),
    .B(net31),
    .C(net37),
    .D(net36),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(net29),
    .B(net38),
    .Y(_01421_));
 sky130_fd_sc_hd__a22oi_2 _07543_ (.A1(net30),
    .A2(net37),
    .B1(net36),
    .B2(net31),
    .Y(_01422_));
 sky130_fd_sc_hd__o21ai_1 _07544_ (.A1(_01421_),
    .A2(_01422_),
    .B1(_01420_),
    .Y(_01423_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(_01244_),
    .A2(_01245_),
    .B1(_01246_),
    .Y(_01424_));
 sky130_fd_sc_hd__a22o_1 _07546_ (.A1(net27),
    .A2(net41),
    .B1(_01244_),
    .B2(_01245_),
    .X(_01425_));
 sky130_fd_sc_hd__a21oi_1 _07547_ (.A1(_01248_),
    .A2(_01425_),
    .B1(_01423_),
    .Y(_01426_));
 sky130_fd_sc_hd__o21bai_2 _07548_ (.A1(_01247_),
    .A2(_01424_),
    .B1_N(_01423_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand3_2 _07549_ (.A(_01248_),
    .B(_01423_),
    .C(_01425_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _07550_ (.A(net27),
    .B(net40),
    .Y(_01429_));
 sky130_fd_sc_hd__a22oi_4 _07551_ (.A1(net28),
    .A2(net39),
    .B1(net40),
    .B2(net27),
    .Y(_01431_));
 sky130_fd_sc_hd__and4_1 _07552_ (.A(net28),
    .B(net27),
    .C(net39),
    .D(net40),
    .X(_01432_));
 sky130_fd_sc_hd__nand4_2 _07553_ (.A(net28),
    .B(net27),
    .C(net39),
    .D(net40),
    .Y(_01433_));
 sky130_fd_sc_hd__o31a_2 _07554_ (.A1(_00044_),
    .A2(_00451_),
    .A3(_01431_),
    .B1(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__o21ai_2 _07555_ (.A1(_01434_),
    .A2(_01426_),
    .B1(_01428_),
    .Y(_01435_));
 sky130_fd_sc_hd__o21a_1 _07556_ (.A1(_01434_),
    .A2(_01426_),
    .B1(_01428_),
    .X(_01436_));
 sky130_fd_sc_hd__o21ai_4 _07557_ (.A1(_01253_),
    .A2(_01416_),
    .B1(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__o211ai_4 _07558_ (.A1(_01239_),
    .A2(_01252_),
    .B1(_01435_),
    .C1(_01417_),
    .Y(_01438_));
 sky130_fd_sc_hd__a22o_1 _07559_ (.A1(net23),
    .A2(net45),
    .B1(_01262_),
    .B2(_01263_),
    .X(_01439_));
 sky130_fd_sc_hd__nand4_2 _07560_ (.A(net26),
    .B(net23),
    .C(net43),
    .D(net42),
    .Y(_01440_));
 sky130_fd_sc_hd__a22o_1 _07561_ (.A1(net23),
    .A2(net43),
    .B1(net42),
    .B2(net26),
    .X(_01442_));
 sky130_fd_sc_hd__nand4_4 _07562_ (.A(_01442_),
    .B(net45),
    .C(net12),
    .D(_01440_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_01440_),
    .B(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__a21o_1 _07564_ (.A1(_01264_),
    .A2(_01439_),
    .B1(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__nand3_1 _07565_ (.A(_01264_),
    .B(_01439_),
    .C(_01444_),
    .Y(_01446_));
 sky130_fd_sc_hd__and4_2 _07566_ (.A(net12),
    .B(net1),
    .C(net46),
    .D(net47),
    .X(_01447_));
 sky130_fd_sc_hd__a22oi_2 _07567_ (.A1(net12),
    .A2(net46),
    .B1(net47),
    .B2(net1),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _07568_ (.A(_01447_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__and3_1 _07569_ (.A(_01445_),
    .B(_01446_),
    .C(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__o2bb2a_1 _07570_ (.A1_N(_01445_),
    .A2_N(_01446_),
    .B1(_01447_),
    .B2(_01448_),
    .X(_01451_));
 sky130_fd_sc_hd__a211oi_1 _07571_ (.A1(_01445_),
    .A2(_01446_),
    .B1(_01447_),
    .C1(_01448_),
    .Y(_01453_));
 sky130_fd_sc_hd__o211a_1 _07572_ (.A1(_01447_),
    .A2(_01448_),
    .B1(_01445_),
    .C1(_01446_),
    .X(_01454_));
 sky130_fd_sc_hd__nor2_1 _07573_ (.A(_01450_),
    .B(_01451_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21bo_1 _07574_ (.A1(_01455_),
    .A2(_01437_),
    .B1_N(_01438_),
    .X(_01456_));
 sky130_fd_sc_hd__a21boi_1 _07575_ (.A1(_01455_),
    .A2(_01437_),
    .B1_N(_01438_),
    .Y(_01457_));
 sky130_fd_sc_hd__a21oi_2 _07576_ (.A1(_01414_),
    .A2(_01415_),
    .B1(_01456_),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_1 _07577_ (.A(_01414_),
    .B(_01456_),
    .Y(_01459_));
 sky130_fd_sc_hd__and3_2 _07578_ (.A(_01414_),
    .B(_01415_),
    .C(_01456_),
    .X(_01460_));
 sky130_fd_sc_hd__nor2_1 _07579_ (.A(_01458_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__o21ai_1 _07580_ (.A1(_01458_),
    .A2(_01460_),
    .B1(_01410_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(_01407_),
    .B(_01461_),
    .Y(_01464_));
 sky130_fd_sc_hd__a21oi_1 _07582_ (.A1(_01407_),
    .A2(_01461_),
    .B1(_01409_),
    .Y(_01465_));
 sky130_fd_sc_hd__o2bb2ai_1 _07583_ (.A1_N(_01224_),
    .A2_N(_01226_),
    .B1(_01280_),
    .B2(_01282_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand4_2 _07584_ (.A(_01224_),
    .B(_01226_),
    .C(_01281_),
    .D(_01283_),
    .Y(_01467_));
 sky130_fd_sc_hd__a21o_1 _07585_ (.A1(_01224_),
    .A2(_01226_),
    .B1(_01284_),
    .X(_01468_));
 sky130_fd_sc_hd__o211ai_2 _07586_ (.A1(_01280_),
    .A2(_01282_),
    .B1(_01224_),
    .C1(_01226_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand3_2 _07587_ (.A(_01465_),
    .B(_01468_),
    .C(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand4_4 _07588_ (.A(_01407_),
    .B(_01462_),
    .C(_01466_),
    .D(_01467_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(_01259_),
    .B(_01261_),
    .Y(_01472_));
 sky130_fd_sc_hd__a22oi_2 _07590_ (.A1(_01268_),
    .A2(_01269_),
    .B1(_01415_),
    .B2(_01459_),
    .Y(_01473_));
 sky130_fd_sc_hd__o2111a_1 _07591_ (.A1(_01457_),
    .A2(_01413_),
    .B1(_01269_),
    .C1(_01268_),
    .D1(_01415_),
    .X(_01475_));
 sky130_fd_sc_hd__nor2_1 _07592_ (.A(_01473_),
    .B(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__a211oi_1 _07593_ (.A1(_01259_),
    .A2(_01261_),
    .B1(_01473_),
    .C1(_01475_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _07594_ (.A(_01472_),
    .B(_01476_),
    .Y(_01478_));
 sky130_fd_sc_hd__o2bb2a_1 _07595_ (.A1_N(_01259_),
    .A2_N(_01261_),
    .B1(_01473_),
    .B2(_01475_),
    .X(_01479_));
 sky130_fd_sc_hd__and3_1 _07596_ (.A(_01476_),
    .B(_01261_),
    .C(_01259_),
    .X(_01480_));
 sky130_fd_sc_hd__nor2_1 _07597_ (.A(_01479_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__a32oi_2 _07598_ (.A1(_01465_),
    .A2(_01468_),
    .A3(_01469_),
    .B1(_01471_),
    .B2(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand3_1 _07599_ (.A(_01299_),
    .B(_01292_),
    .C(_01291_),
    .Y(_01483_));
 sky130_fd_sc_hd__a21o_1 _07600_ (.A1(_01291_),
    .A2(_01292_),
    .B1(_01299_),
    .X(_01484_));
 sky130_fd_sc_hd__a21oi_1 _07601_ (.A1(_01483_),
    .A2(_01484_),
    .B1(_01482_),
    .Y(_01486_));
 sky130_fd_sc_hd__nand3_1 _07602_ (.A(_01482_),
    .B(_01483_),
    .C(_01484_),
    .Y(_01487_));
 sky130_fd_sc_hd__a21o_1 _07603_ (.A1(_01476_),
    .A2(_01472_),
    .B1(_01473_),
    .X(_01488_));
 sky130_fd_sc_hd__inv_2 _07604_ (.A(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__o21a_2 _07605_ (.A1(_01486_),
    .A2(_01489_),
    .B1(_01487_),
    .X(_01490_));
 sky130_fd_sc_hd__and2b_1 _07606_ (.A_N(_01490_),
    .B(_01312_),
    .X(_01491_));
 sky130_fd_sc_hd__inv_2 _07607_ (.A(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__xnor2_4 _07608_ (.A(_01312_),
    .B(_01490_),
    .Y(_01493_));
 sky130_fd_sc_hd__o2bb2ai_4 _07609_ (.A1_N(_01407_),
    .A2_N(_01410_),
    .B1(_01458_),
    .B2(_01460_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand3_2 _07610_ (.A(_01407_),
    .B(_01410_),
    .C(_01461_),
    .Y(_01495_));
 sky130_fd_sc_hd__o211ai_1 _07611_ (.A1(_01458_),
    .A2(_01460_),
    .B1(_01407_),
    .C1(_01410_),
    .Y(_01497_));
 sky130_fd_sc_hd__a21bo_1 _07612_ (.A1(_01407_),
    .A2(_01410_),
    .B1_N(_01461_),
    .X(_01498_));
 sky130_fd_sc_hd__o22ai_4 _07613_ (.A1(_01394_),
    .A2(_01395_),
    .B1(_01398_),
    .B2(_01370_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(net9),
    .B(net33),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_2 _07615_ (.A(net9),
    .B(net44),
    .Y(_01501_));
 sky130_fd_sc_hd__nand4_2 _07616_ (.A(net9),
    .B(net10),
    .C(net44),
    .D(net33),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _07617_ (.A(net8),
    .B(net55),
    .Y(_01503_));
 sky130_fd_sc_hd__a22oi_1 _07618_ (.A1(net9),
    .A2(net44),
    .B1(net33),
    .B2(net10),
    .Y(_01504_));
 sky130_fd_sc_hd__nand3_1 _07619_ (.A(_01501_),
    .B(net33),
    .C(net10),
    .Y(_01505_));
 sky130_fd_sc_hd__nand3_1 _07620_ (.A(_01314_),
    .B(net44),
    .C(net9),
    .Y(_01506_));
 sky130_fd_sc_hd__nand4b_4 _07621_ (.A_N(_01504_),
    .B(net55),
    .C(net8),
    .D(_01502_),
    .Y(_01508_));
 sky130_fd_sc_hd__o21ai_1 _07622_ (.A1(_01503_),
    .A2(_01504_),
    .B1(_01502_),
    .Y(_01509_));
 sky130_fd_sc_hd__o211ai_2 _07623_ (.A1(_00198_),
    .A2(_00341_),
    .B1(_01319_),
    .C1(_01321_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand3_2 _07624_ (.A(_01322_),
    .B(_01509_),
    .C(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__a21o_1 _07625_ (.A1(_01322_),
    .A2(_01510_),
    .B1(_01509_),
    .X(_01512_));
 sky130_fd_sc_hd__a22oi_4 _07626_ (.A1(net8),
    .A2(net58),
    .B1(net59),
    .B2(net7),
    .Y(_01513_));
 sky130_fd_sc_hd__a22o_1 _07627_ (.A1(net8),
    .A2(net58),
    .B1(net59),
    .B2(net7),
    .X(_01514_));
 sky130_fd_sc_hd__and4_1 _07628_ (.A(net7),
    .B(net8),
    .C(net58),
    .D(net59),
    .X(_01515_));
 sky130_fd_sc_hd__nand4_1 _07629_ (.A(net7),
    .B(net8),
    .C(net58),
    .D(net59),
    .Y(_01516_));
 sky130_fd_sc_hd__a211o_1 _07630_ (.A1(net6),
    .A2(net60),
    .B1(_01513_),
    .C1(_01515_),
    .X(_01517_));
 sky130_fd_sc_hd__o211ai_1 _07631_ (.A1(_01513_),
    .A2(_01515_),
    .B1(net6),
    .C1(net60),
    .Y(_01519_));
 sky130_fd_sc_hd__o22a_1 _07632_ (.A1(_00187_),
    .A2(_00352_),
    .B1(_01513_),
    .B2(_01515_),
    .X(_01520_));
 sky130_fd_sc_hd__and4_1 _07633_ (.A(_01514_),
    .B(_01516_),
    .C(net6),
    .D(net60),
    .X(_01521_));
 sky130_fd_sc_hd__nand2_1 _07634_ (.A(_01517_),
    .B(_01519_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand3_2 _07635_ (.A(_01511_),
    .B(_01512_),
    .C(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__a21boi_2 _07636_ (.A1(_01512_),
    .A2(_01522_),
    .B1_N(_01511_),
    .Y(_01524_));
 sky130_fd_sc_hd__a21bo_1 _07637_ (.A1(_01512_),
    .A2(_01522_),
    .B1_N(_01511_),
    .X(_01525_));
 sky130_fd_sc_hd__a21oi_2 _07638_ (.A1(_01327_),
    .A2(_01328_),
    .B1(_01341_),
    .Y(_01526_));
 sky130_fd_sc_hd__o2bb2ai_2 _07639_ (.A1_N(_01327_),
    .A2_N(_01328_),
    .B1(_01335_),
    .B2(_01336_),
    .Y(_01527_));
 sky130_fd_sc_hd__a21oi_2 _07640_ (.A1(_01344_),
    .A2(_01527_),
    .B1(_01525_),
    .Y(_01528_));
 sky130_fd_sc_hd__o21ai_2 _07641_ (.A1(_01343_),
    .A2(_01526_),
    .B1(_01524_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor3_1 _07642_ (.A(_01343_),
    .B(_01524_),
    .C(_01526_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand3_4 _07643_ (.A(_01344_),
    .B(_01525_),
    .C(_01527_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(net4),
    .B(net61),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _07645_ (.A(net4),
    .B(net62),
    .Y(_01534_));
 sky130_fd_sc_hd__and4_2 _07646_ (.A(net5),
    .B(net4),
    .C(net62),
    .D(net61),
    .X(_01535_));
 sky130_fd_sc_hd__nand4_1 _07647_ (.A(net5),
    .B(net4),
    .C(net62),
    .D(net61),
    .Y(_01536_));
 sky130_fd_sc_hd__a22o_1 _07648_ (.A1(net4),
    .A2(net62),
    .B1(net61),
    .B2(net5),
    .X(_01537_));
 sky130_fd_sc_hd__nand3_1 _07649_ (.A(_01534_),
    .B(net61),
    .C(net5),
    .Y(_01538_));
 sky130_fd_sc_hd__nand3_1 _07650_ (.A(_01360_),
    .B(net62),
    .C(net4),
    .Y(_01539_));
 sky130_fd_sc_hd__and4_2 _07651_ (.A(_01537_),
    .B(net63),
    .C(net3),
    .D(_01536_),
    .X(_01541_));
 sky130_fd_sc_hd__nand4_2 _07652_ (.A(_01537_),
    .B(net63),
    .C(net3),
    .D(_01536_),
    .Y(_01542_));
 sky130_fd_sc_hd__o21a_1 _07653_ (.A1(_00187_),
    .A2(_00352_),
    .B1(_01516_),
    .X(_01543_));
 sky130_fd_sc_hd__a31o_1 _07654_ (.A1(_01514_),
    .A2(net60),
    .A3(net6),
    .B1(_01515_),
    .X(_01544_));
 sky130_fd_sc_hd__a22oi_4 _07655_ (.A1(net4),
    .A2(net63),
    .B1(_01359_),
    .B2(_01361_),
    .Y(_01545_));
 sky130_fd_sc_hd__and4_2 _07656_ (.A(_01359_),
    .B(_01361_),
    .C(net4),
    .D(net63),
    .X(_01546_));
 sky130_fd_sc_hd__nand4_1 _07657_ (.A(_01359_),
    .B(_01361_),
    .C(net4),
    .D(net63),
    .Y(_01547_));
 sky130_fd_sc_hd__o22ai_4 _07658_ (.A1(_01513_),
    .A2(_01543_),
    .B1(_01545_),
    .B2(_01546_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand3b_2 _07659_ (.A_N(_01545_),
    .B(_01547_),
    .C(_01544_),
    .Y(_01549_));
 sky130_fd_sc_hd__o211a_1 _07660_ (.A1(_01535_),
    .A2(_01541_),
    .B1(_01548_),
    .C1(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__o211ai_4 _07661_ (.A1(_01535_),
    .A2(_01541_),
    .B1(_01548_),
    .C1(_01549_),
    .Y(_01552_));
 sky130_fd_sc_hd__a211oi_2 _07662_ (.A1(_01548_),
    .A2(_01549_),
    .B1(_01535_),
    .C1(_01541_),
    .Y(_01553_));
 sky130_fd_sc_hd__a211o_1 _07663_ (.A1(_01548_),
    .A2(_01549_),
    .B1(_01535_),
    .C1(_01541_),
    .X(_01554_));
 sky130_fd_sc_hd__nor2_1 _07664_ (.A(_01550_),
    .B(_01553_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(_01552_),
    .B(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__o32a_1 _07666_ (.A1(_01343_),
    .A2(_01524_),
    .A3(_01526_),
    .B1(_01550_),
    .B2(_01553_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _07667_ (.A(_01555_),
    .B(_01530_),
    .Y(_01558_));
 sky130_fd_sc_hd__o21ai_1 _07668_ (.A1(_01528_),
    .A2(_01556_),
    .B1(_01532_),
    .Y(_01559_));
 sky130_fd_sc_hd__nand3b_2 _07669_ (.A_N(_01349_),
    .B(_01351_),
    .C(_01367_),
    .Y(_01560_));
 sky130_fd_sc_hd__o21bai_2 _07670_ (.A1(_01349_),
    .A2(_01350_),
    .B1_N(_01367_),
    .Y(_01561_));
 sky130_fd_sc_hd__o21ai_1 _07671_ (.A1(_01349_),
    .A2(_01350_),
    .B1(_01367_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand4b_1 _07672_ (.A_N(_01349_),
    .B(_01351_),
    .C(_01365_),
    .D(_01366_),
    .Y(_01564_));
 sky130_fd_sc_hd__o211ai_4 _07673_ (.A1(_01528_),
    .A2(_01557_),
    .B1(_01560_),
    .C1(_01561_),
    .Y(_01565_));
 sky130_fd_sc_hd__inv_2 _07674_ (.A(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__a22oi_2 _07675_ (.A1(_01532_),
    .A2(_01558_),
    .B1(_01560_),
    .B2(_01561_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand3_2 _07676_ (.A(_01559_),
    .B(_01563_),
    .C(_01564_),
    .Y(_01568_));
 sky130_fd_sc_hd__o41ai_4 _07677_ (.A1(_01513_),
    .A2(_01543_),
    .A3(_01545_),
    .A4(_01546_),
    .B1(_01552_),
    .Y(_01569_));
 sky130_fd_sc_hd__o2bb2ai_2 _07678_ (.A1_N(_01389_),
    .A2_N(_01390_),
    .B1(_01391_),
    .B2(_01233_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand4_4 _07679_ (.A(_01234_),
    .B(_01389_),
    .C(_01390_),
    .D(_01392_),
    .Y(_01571_));
 sky130_fd_sc_hd__a21oi_2 _07680_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01569_),
    .Y(_01572_));
 sky130_fd_sc_hd__a21o_1 _07681_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01569_),
    .X(_01574_));
 sky130_fd_sc_hd__nand3_4 _07682_ (.A(_01569_),
    .B(_01570_),
    .C(_01571_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(net32),
    .B(net64),
    .Y(_01576_));
 sky130_fd_sc_hd__nand2_1 _07684_ (.A(net32),
    .B(net34),
    .Y(_01577_));
 sky130_fd_sc_hd__and2_1 _07685_ (.A(net31),
    .B(net35),
    .X(_01578_));
 sky130_fd_sc_hd__a22o_1 _07686_ (.A1(net2),
    .A2(net64),
    .B1(net34),
    .B2(net32),
    .X(_01579_));
 sky130_fd_sc_hd__nand3_1 _07687_ (.A(_01577_),
    .B(net64),
    .C(net2),
    .Y(_01580_));
 sky130_fd_sc_hd__nand3_1 _07688_ (.A(_01378_),
    .B(net34),
    .C(net32),
    .Y(_01581_));
 sky130_fd_sc_hd__o2111ai_4 _07689_ (.A1(_01379_),
    .A2(_01576_),
    .B1(net31),
    .C1(net35),
    .D1(_01579_),
    .Y(_01582_));
 sky130_fd_sc_hd__o2bb2ai_2 _07690_ (.A1_N(_01578_),
    .A2_N(_01579_),
    .B1(_01379_),
    .B2(_01576_),
    .Y(_01583_));
 sky130_fd_sc_hd__o211a_1 _07691_ (.A1(_00110_),
    .A2(_00407_),
    .B1(_01382_),
    .C1(_01383_),
    .X(_01585_));
 sky130_fd_sc_hd__o211ai_2 _07692_ (.A1(_00110_),
    .A2(_00407_),
    .B1(_01382_),
    .C1(_01383_),
    .Y(_01586_));
 sky130_fd_sc_hd__a21oi_1 _07693_ (.A1(_01384_),
    .A2(_01586_),
    .B1(_01583_),
    .Y(_01587_));
 sky130_fd_sc_hd__a21o_1 _07694_ (.A1(_01384_),
    .A2(_01586_),
    .B1(_01583_),
    .X(_01588_));
 sky130_fd_sc_hd__nand2_1 _07695_ (.A(_01384_),
    .B(_01583_),
    .Y(_01589_));
 sky130_fd_sc_hd__and3_1 _07696_ (.A(_01384_),
    .B(_01583_),
    .C(_01586_),
    .X(_01590_));
 sky130_fd_sc_hd__a211o_1 _07697_ (.A1(net29),
    .A2(net38),
    .B1(_01418_),
    .C1(_01422_),
    .X(_01591_));
 sky130_fd_sc_hd__o211ai_2 _07698_ (.A1(_01418_),
    .A2(_01422_),
    .B1(net29),
    .C1(net38),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_01591_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__a2bb2o_1 _07700_ (.A1_N(_01585_),
    .A2_N(_01589_),
    .B1(_01588_),
    .B2(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__o2bb2a_1 _07701_ (.A1_N(_01593_),
    .A2_N(_01588_),
    .B1(_01585_),
    .B2(_01589_),
    .X(_01596_));
 sky130_fd_sc_hd__a21oi_2 _07702_ (.A1(_01574_),
    .A2(_01575_),
    .B1(_01594_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21o_1 _07703_ (.A1(_01574_),
    .A2(_01575_),
    .B1(_01594_),
    .X(_01598_));
 sky130_fd_sc_hd__and3_1 _07704_ (.A(_01574_),
    .B(_01575_),
    .C(_01594_),
    .X(_01599_));
 sky130_fd_sc_hd__nand3_1 _07705_ (.A(_01574_),
    .B(_01575_),
    .C(_01594_),
    .Y(_01600_));
 sky130_fd_sc_hd__o21a_1 _07706_ (.A1(_01597_),
    .A2(_01599_),
    .B1(_01568_),
    .X(_01601_));
 sky130_fd_sc_hd__nand3_1 _07707_ (.A(_01565_),
    .B(_01598_),
    .C(_01600_),
    .Y(_01602_));
 sky130_fd_sc_hd__a31o_1 _07708_ (.A1(_01565_),
    .A2(_01598_),
    .A3(_01600_),
    .B1(_01567_),
    .X(_01603_));
 sky130_fd_sc_hd__o2bb2ai_2 _07709_ (.A1_N(_01400_),
    .A2_N(_01499_),
    .B1(_01566_),
    .B2(_01601_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand3_4 _07710_ (.A(_01603_),
    .B(_01499_),
    .C(_01400_),
    .Y(_01605_));
 sky130_fd_sc_hd__o21ai_1 _07711_ (.A1(_01596_),
    .A2(_01572_),
    .B1(_01575_),
    .Y(_01607_));
 sky130_fd_sc_hd__o211ai_2 _07712_ (.A1(_01450_),
    .A2(_01451_),
    .B1(_01437_),
    .C1(_01438_),
    .Y(_01608_));
 sky130_fd_sc_hd__o2bb2ai_1 _07713_ (.A1_N(_01437_),
    .A2_N(_01438_),
    .B1(_01453_),
    .B2(_01454_),
    .Y(_01609_));
 sky130_fd_sc_hd__o211ai_1 _07714_ (.A1(_01453_),
    .A2(_01454_),
    .B1(_01437_),
    .C1(_01438_),
    .Y(_01610_));
 sky130_fd_sc_hd__o2bb2ai_1 _07715_ (.A1_N(_01437_),
    .A2_N(_01438_),
    .B1(_01450_),
    .B2(_01451_),
    .Y(_01611_));
 sky130_fd_sc_hd__o2111ai_4 _07716_ (.A1(_01596_),
    .A2(_01572_),
    .B1(_01575_),
    .C1(_01608_),
    .D1(_01609_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand3_2 _07717_ (.A(_01611_),
    .B(_01607_),
    .C(_01610_),
    .Y(_01613_));
 sky130_fd_sc_hd__a22oi_4 _07718_ (.A1(net29),
    .A2(net37),
    .B1(net36),
    .B2(net30),
    .Y(_01614_));
 sky130_fd_sc_hd__and4_2 _07719_ (.A(net30),
    .B(net29),
    .C(net37),
    .D(net36),
    .X(_01615_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(net28),
    .B(net38),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _07721_ (.A(_01616_),
    .B(_01614_),
    .Y(_01618_));
 sky130_fd_sc_hd__o21bai_1 _07722_ (.A1(_01614_),
    .A2(_01616_),
    .B1_N(_01615_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand4b_4 _07723_ (.A_N(_01431_),
    .B(_01433_),
    .C(net26),
    .D(net41),
    .Y(_01620_));
 sky130_fd_sc_hd__o22ai_4 _07724_ (.A1(_00044_),
    .A2(_00451_),
    .B1(_01431_),
    .B2(_01432_),
    .Y(_01621_));
 sky130_fd_sc_hd__o211a_2 _07725_ (.A1(_01615_),
    .A2(_01618_),
    .B1(_01620_),
    .C1(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__o211ai_4 _07726_ (.A1(_01615_),
    .A2(_01618_),
    .B1(_01620_),
    .C1(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(net26),
    .B(net39),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_2 _07728_ (.A(net26),
    .B(net40),
    .Y(_01625_));
 sky130_fd_sc_hd__and4_1 _07729_ (.A(net26),
    .B(net27),
    .C(net39),
    .D(net40),
    .X(_01626_));
 sky130_fd_sc_hd__nand4_2 _07730_ (.A(net26),
    .B(net27),
    .C(net39),
    .D(net40),
    .Y(_01627_));
 sky130_fd_sc_hd__a22o_2 _07731_ (.A1(net27),
    .A2(net39),
    .B1(net40),
    .B2(net26),
    .X(_01629_));
 sky130_fd_sc_hd__o2111a_2 _07732_ (.A1(_01429_),
    .A2(_01624_),
    .B1(net23),
    .C1(net41),
    .D1(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__o2111ai_4 _07733_ (.A1(_01429_),
    .A2(_01624_),
    .B1(net23),
    .C1(net41),
    .D1(_01629_),
    .Y(_01631_));
 sky130_fd_sc_hd__o31a_1 _07734_ (.A1(_00077_),
    .A2(_00440_),
    .A3(_01625_),
    .B1(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__a21oi_2 _07735_ (.A1(_01620_),
    .A2(_01621_),
    .B1(_01619_),
    .Y(_01633_));
 sky130_fd_sc_hd__a21o_1 _07736_ (.A1(_01620_),
    .A2(_01621_),
    .B1(_01619_),
    .X(_01634_));
 sky130_fd_sc_hd__o21ai_2 _07737_ (.A1(_01626_),
    .A2(_01630_),
    .B1(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__o211ai_4 _07738_ (.A1(_01626_),
    .A2(_01630_),
    .B1(_01634_),
    .C1(_01623_),
    .Y(_01636_));
 sky130_fd_sc_hd__o21ai_1 _07739_ (.A1(_01632_),
    .A2(_01633_),
    .B1(_01623_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21o_1 _07740_ (.A1(_01427_),
    .A2(_01428_),
    .B1(_01434_),
    .X(_01638_));
 sky130_fd_sc_hd__nand3_1 _07741_ (.A(_01427_),
    .B(_01428_),
    .C(_01434_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand3b_1 _07742_ (.A_N(_01434_),
    .B(_01428_),
    .C(_01427_),
    .Y(_01641_));
 sky130_fd_sc_hd__a21bo_1 _07743_ (.A1(_01427_),
    .A2(_01428_),
    .B1_N(_01434_),
    .X(_01642_));
 sky130_fd_sc_hd__nand4_2 _07744_ (.A(_01623_),
    .B(_01636_),
    .C(_01638_),
    .D(_01640_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand3_2 _07745_ (.A(_01637_),
    .B(_01641_),
    .C(_01642_),
    .Y(_01644_));
 sky130_fd_sc_hd__and4_1 _07746_ (.A(net12),
    .B(net23),
    .C(net43),
    .D(net42),
    .X(_01645_));
 sky130_fd_sc_hd__nand4_1 _07747_ (.A(net12),
    .B(net23),
    .C(net43),
    .D(net42),
    .Y(_01646_));
 sky130_fd_sc_hd__a22o_1 _07748_ (.A1(net12),
    .A2(net43),
    .B1(net42),
    .B2(net23),
    .X(_01647_));
 sky130_fd_sc_hd__and4_2 _07749_ (.A(_01647_),
    .B(net45),
    .C(net1),
    .D(_01646_),
    .X(_01648_));
 sky130_fd_sc_hd__a31o_1 _07750_ (.A1(_01647_),
    .A2(net45),
    .A3(net1),
    .B1(_01645_),
    .X(_01649_));
 sky130_fd_sc_hd__a22o_1 _07751_ (.A1(net12),
    .A2(net45),
    .B1(_01440_),
    .B2(_01442_),
    .X(_01651_));
 sky130_fd_sc_hd__a21o_1 _07752_ (.A1(_01443_),
    .A2(_01651_),
    .B1(_01649_),
    .X(_01652_));
 sky130_fd_sc_hd__o211ai_4 _07753_ (.A1(_01645_),
    .A2(_01648_),
    .B1(_01651_),
    .C1(_01443_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__and4_1 _07755_ (.A(_01652_),
    .B(_01653_),
    .C(net1),
    .D(net46),
    .X(_01655_));
 sky130_fd_sc_hd__o2bb2a_1 _07756_ (.A1_N(_01652_),
    .A2_N(_01653_),
    .B1(_00033_),
    .B2(_00484_),
    .X(_01656_));
 sky130_fd_sc_hd__a211o_1 _07757_ (.A1(_01652_),
    .A2(_01653_),
    .B1(_00033_),
    .C1(_00484_),
    .X(_01657_));
 sky130_fd_sc_hd__o211ai_2 _07758_ (.A1(_00033_),
    .A2(_00484_),
    .B1(_01652_),
    .C1(_01653_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _07759_ (.A(_01657_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__a21bo_1 _07760_ (.A1(_01659_),
    .A2(_01643_),
    .B1_N(_01644_),
    .X(_01660_));
 sky130_fd_sc_hd__nand3_2 _07761_ (.A(_01612_),
    .B(_01613_),
    .C(_01660_),
    .Y(_01662_));
 sky130_fd_sc_hd__inv_2 _07762_ (.A(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21o_1 _07763_ (.A1(_01612_),
    .A2(_01613_),
    .B1(_01660_),
    .X(_01664_));
 sky130_fd_sc_hd__inv_2 _07764_ (.A(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(_01662_),
    .B(_01664_),
    .Y(_01666_));
 sky130_fd_sc_hd__nand3_1 _07766_ (.A(_01604_),
    .B(_01662_),
    .C(_01664_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_4 _07767_ (.A(_01605_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__inv_2 _07768_ (.A(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__a21oi_4 _07769_ (.A1(_01494_),
    .A2(_01495_),
    .B1(_01668_),
    .Y(_01670_));
 sky130_fd_sc_hd__a21o_1 _07770_ (.A1(_01494_),
    .A2(_01495_),
    .B1(_01668_),
    .X(_01671_));
 sky130_fd_sc_hd__o211a_1 _07771_ (.A1(_01409_),
    .A2(_01464_),
    .B1(_01668_),
    .C1(_01494_),
    .X(_01673_));
 sky130_fd_sc_hd__o211ai_2 _07772_ (.A1(_01409_),
    .A2(_01464_),
    .B1(_01668_),
    .C1(_01494_),
    .Y(_01674_));
 sky130_fd_sc_hd__a31o_1 _07773_ (.A1(_01264_),
    .A2(_01439_),
    .A3(_01444_),
    .B1(_01450_),
    .X(_01675_));
 sky130_fd_sc_hd__a21boi_1 _07774_ (.A1(_01612_),
    .A2(_01660_),
    .B1_N(_01613_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21boi_2 _07775_ (.A1(_01613_),
    .A2(_01662_),
    .B1_N(_01675_),
    .Y(_01677_));
 sky130_fd_sc_hd__xnor2_2 _07776_ (.A(_01675_),
    .B(_01676_),
    .Y(_01678_));
 sky130_fd_sc_hd__and2_1 _07777_ (.A(_01447_),
    .B(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__xor2_1 _07778_ (.A(_01447_),
    .B(_01678_),
    .X(_01680_));
 sky130_fd_sc_hd__xnor2_2 _07779_ (.A(_01447_),
    .B(_01678_),
    .Y(_01681_));
 sky130_fd_sc_hd__a31oi_2 _07780_ (.A1(_01494_),
    .A2(_01495_),
    .A3(_01668_),
    .B1(_01680_),
    .Y(_01682_));
 sky130_fd_sc_hd__a32oi_2 _07781_ (.A1(_01497_),
    .A2(_01498_),
    .A3(_01669_),
    .B1(_01674_),
    .B2(_01681_),
    .Y(_01684_));
 sky130_fd_sc_hd__o2bb2ai_2 _07782_ (.A1_N(_01470_),
    .A2_N(_01471_),
    .B1(_01479_),
    .B2(_01480_),
    .Y(_01685_));
 sky130_fd_sc_hd__o211ai_2 _07783_ (.A1(_01477_),
    .A2(_01478_),
    .B1(_01470_),
    .C1(_01471_),
    .Y(_01686_));
 sky130_fd_sc_hd__o211ai_1 _07784_ (.A1(_01479_),
    .A2(_01480_),
    .B1(_01470_),
    .C1(_01471_),
    .Y(_01687_));
 sky130_fd_sc_hd__o2bb2ai_1 _07785_ (.A1_N(_01470_),
    .A2_N(_01471_),
    .B1(_01477_),
    .B2(_01478_),
    .Y(_01688_));
 sky130_fd_sc_hd__a2bb2oi_1 _07786_ (.A1_N(_01670_),
    .A2_N(_01682_),
    .B1(_01687_),
    .B2(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__o211ai_4 _07787_ (.A1(_01670_),
    .A2(_01682_),
    .B1(_01685_),
    .C1(_01686_),
    .Y(_01690_));
 sky130_fd_sc_hd__a21boi_1 _07788_ (.A1(_01685_),
    .A2(_01686_),
    .B1_N(_01684_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand3_1 _07789_ (.A(_01688_),
    .B(_01684_),
    .C(_01687_),
    .Y(_01692_));
 sky130_fd_sc_hd__a21oi_1 _07790_ (.A1(_01447_),
    .A2(_01678_),
    .B1(_01677_),
    .Y(_01693_));
 sky130_fd_sc_hd__or3_2 _07791_ (.A(_01677_),
    .B(_01679_),
    .C(_01691_),
    .X(_01695_));
 sky130_fd_sc_hd__nand2b_1 _07792_ (.A_N(_01486_),
    .B(_01487_),
    .Y(_01696_));
 sky130_fd_sc_hd__or2_1 _07793_ (.A(_01489_),
    .B(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__inv_2 _07794_ (.A(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(_01696_),
    .B(_01489_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand3_2 _07796_ (.A(_01690_),
    .B(_01695_),
    .C(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__o2bb2ai_2 _07797_ (.A1_N(_01511_),
    .A2_N(_01512_),
    .B1(_01520_),
    .B2(_01521_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_2 _07798_ (.A(_01523_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_2 _07799_ (.A(net8),
    .B(net33),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_2 _07800_ (.A(net8),
    .B(net44),
    .Y(_01704_));
 sky130_fd_sc_hd__and4_1 _07801_ (.A(net9),
    .B(net8),
    .C(net44),
    .D(net33),
    .X(_01706_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(net7),
    .B(net55),
    .Y(_01707_));
 sky130_fd_sc_hd__a22oi_4 _07803_ (.A1(net8),
    .A2(net44),
    .B1(net33),
    .B2(net9),
    .Y(_01708_));
 sky130_fd_sc_hd__a22o_1 _07804_ (.A1(net8),
    .A2(net44),
    .B1(net33),
    .B2(net9),
    .X(_01709_));
 sky130_fd_sc_hd__nand3_1 _07805_ (.A(_01704_),
    .B(net33),
    .C(net9),
    .Y(_01710_));
 sky130_fd_sc_hd__nand3_1 _07806_ (.A(_01500_),
    .B(net44),
    .C(net8),
    .Y(_01711_));
 sky130_fd_sc_hd__o2111ai_4 _07807_ (.A1(_01501_),
    .A2(_01703_),
    .B1(net7),
    .C1(net55),
    .D1(_01709_),
    .Y(_01712_));
 sky130_fd_sc_hd__o22ai_4 _07808_ (.A1(_01501_),
    .A2(_01703_),
    .B1(_01707_),
    .B2(_01708_),
    .Y(_01713_));
 sky130_fd_sc_hd__o211ai_4 _07809_ (.A1(_00209_),
    .A2(_00341_),
    .B1(_01505_),
    .C1(_01506_),
    .Y(_01714_));
 sky130_fd_sc_hd__and3_2 _07810_ (.A(_01508_),
    .B(_01713_),
    .C(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__nand3_2 _07811_ (.A(_01508_),
    .B(_01713_),
    .C(_01714_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(net5),
    .B(net60),
    .Y(_01718_));
 sky130_fd_sc_hd__a22oi_4 _07813_ (.A1(net7),
    .A2(net58),
    .B1(net59),
    .B2(net6),
    .Y(_01719_));
 sky130_fd_sc_hd__and4_1 _07814_ (.A(net7),
    .B(net6),
    .C(net58),
    .D(net59),
    .X(_01720_));
 sky130_fd_sc_hd__nand4_1 _07815_ (.A(net7),
    .B(net6),
    .C(net58),
    .D(net59),
    .Y(_01721_));
 sky130_fd_sc_hd__a211o_1 _07816_ (.A1(net5),
    .A2(net60),
    .B1(_01719_),
    .C1(_01720_),
    .X(_01722_));
 sky130_fd_sc_hd__o211ai_4 _07817_ (.A1(_01719_),
    .A2(_01720_),
    .B1(net5),
    .C1(net60),
    .Y(_01723_));
 sky130_fd_sc_hd__o22a_1 _07818_ (.A1(_00154_),
    .A2(_00352_),
    .B1(_01719_),
    .B2(_01720_),
    .X(_01724_));
 sky130_fd_sc_hd__and4b_1 _07819_ (.A_N(_01719_),
    .B(_01721_),
    .C(net5),
    .D(net60),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_01722_),
    .B(_01723_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21oi_4 _07821_ (.A1(_01508_),
    .A2(_01714_),
    .B1(_01713_),
    .Y(_01728_));
 sky130_fd_sc_hd__a21o_1 _07822_ (.A1(_01508_),
    .A2(_01714_),
    .B1(_01713_),
    .X(_01729_));
 sky130_fd_sc_hd__a21oi_1 _07823_ (.A1(_01722_),
    .A2(_01723_),
    .B1(_01728_),
    .Y(_01730_));
 sky130_fd_sc_hd__and3_1 _07824_ (.A(_01717_),
    .B(_01722_),
    .C(_01723_),
    .X(_01731_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_01717_),
    .B(_01726_),
    .C(_01729_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21oi_2 _07826_ (.A1(_01726_),
    .A2(_01729_),
    .B1(_01715_),
    .Y(_01733_));
 sky130_fd_sc_hd__o211a_2 _07827_ (.A1(_01715_),
    .A2(_01730_),
    .B1(_01523_),
    .C1(_01701_),
    .X(_01734_));
 sky130_fd_sc_hd__o211ai_2 _07828_ (.A1(_01715_),
    .A2(_01730_),
    .B1(_01523_),
    .C1(_01701_),
    .Y(_01735_));
 sky130_fd_sc_hd__o2bb2ai_2 _07829_ (.A1_N(_01523_),
    .A2_N(_01701_),
    .B1(_01728_),
    .B2(_01731_),
    .Y(_01736_));
 sky130_fd_sc_hd__nand2_2 _07830_ (.A(net3),
    .B(net62),
    .Y(_01737_));
 sky130_fd_sc_hd__nand4_4 _07831_ (.A(net3),
    .B(net4),
    .C(net62),
    .D(net61),
    .Y(_01739_));
 sky130_fd_sc_hd__a22o_1 _07832_ (.A1(net3),
    .A2(net62),
    .B1(net61),
    .B2(net4),
    .X(_01740_));
 sky130_fd_sc_hd__nand3_1 _07833_ (.A(_01737_),
    .B(net61),
    .C(net4),
    .Y(_01741_));
 sky130_fd_sc_hd__nand3_1 _07834_ (.A(_01533_),
    .B(net62),
    .C(net3),
    .Y(_01742_));
 sky130_fd_sc_hd__nand4_4 _07835_ (.A(_01740_),
    .B(net63),
    .C(net2),
    .D(_01739_),
    .Y(_01743_));
 sky130_fd_sc_hd__o31a_1 _07836_ (.A1(_00132_),
    .A2(_00374_),
    .A3(_01533_),
    .B1(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__o21ai_1 _07837_ (.A1(_01533_),
    .A2(_01737_),
    .B1(_01743_),
    .Y(_01745_));
 sky130_fd_sc_hd__o211a_1 _07838_ (.A1(_00132_),
    .A2(_00396_),
    .B1(_01538_),
    .C1(_01539_),
    .X(_01746_));
 sky130_fd_sc_hd__o211ai_2 _07839_ (.A1(_00132_),
    .A2(_00396_),
    .B1(_01538_),
    .C1(_01539_),
    .Y(_01747_));
 sky130_fd_sc_hd__o21a_1 _07840_ (.A1(_00154_),
    .A2(_00352_),
    .B1(_01721_),
    .X(_01748_));
 sky130_fd_sc_hd__o21ai_1 _07841_ (.A1(_01718_),
    .A2(_01719_),
    .B1(_01721_),
    .Y(_01750_));
 sky130_fd_sc_hd__o2bb2ai_2 _07842_ (.A1_N(_01542_),
    .A2_N(_01747_),
    .B1(_01748_),
    .B2(_01719_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_01750_),
    .B(_01542_),
    .Y(_01752_));
 sky130_fd_sc_hd__nand3_1 _07844_ (.A(_01750_),
    .B(_01747_),
    .C(_01542_),
    .Y(_01753_));
 sky130_fd_sc_hd__a22oi_2 _07845_ (.A1(_01739_),
    .A2(_01743_),
    .B1(_01751_),
    .B2(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__a22o_1 _07846_ (.A1(_01739_),
    .A2(_01743_),
    .B1(_01751_),
    .B2(_01753_),
    .X(_01755_));
 sky130_fd_sc_hd__o211a_1 _07847_ (.A1(_01746_),
    .A2(_01752_),
    .B1(_01751_),
    .C1(_01744_),
    .X(_01756_));
 sky130_fd_sc_hd__o211ai_1 _07848_ (.A1(_01746_),
    .A2(_01752_),
    .B1(_01751_),
    .C1(_01744_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(_01755_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _07850_ (.A(_01754_),
    .B(_01756_),
    .Y(_01759_));
 sky130_fd_sc_hd__a21oi_2 _07851_ (.A1(_01702_),
    .A2(_01733_),
    .B1(_01759_),
    .Y(_01761_));
 sky130_fd_sc_hd__o21ai_2 _07852_ (.A1(_01754_),
    .A2(_01756_),
    .B1(_01736_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _07853_ (.A(_01735_),
    .B(_01759_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _07854_ (.A(_01736_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__o211ai_2 _07855_ (.A1(_01550_),
    .A2(_01553_),
    .B1(_01530_),
    .C1(_01532_),
    .Y(_01765_));
 sky130_fd_sc_hd__o21ai_1 _07856_ (.A1(_01528_),
    .A2(_01531_),
    .B1(_01555_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand4_2 _07857_ (.A(_01530_),
    .B(_01532_),
    .C(_01552_),
    .D(_01554_),
    .Y(_01767_));
 sky130_fd_sc_hd__o2bb2ai_1 _07858_ (.A1_N(_01530_),
    .A2_N(_01532_),
    .B1(_01550_),
    .B2(_01553_),
    .Y(_01768_));
 sky130_fd_sc_hd__o211ai_4 _07859_ (.A1(_01734_),
    .A2(_01761_),
    .B1(_01767_),
    .C1(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand3_4 _07860_ (.A(_01766_),
    .B(_01764_),
    .C(_01765_),
    .Y(_01770_));
 sky130_fd_sc_hd__a2bb2o_1 _07861_ (.A1_N(_01746_),
    .A2_N(_01752_),
    .B1(_01751_),
    .B2(_01745_),
    .X(_01772_));
 sky130_fd_sc_hd__o2bb2a_1 _07862_ (.A1_N(_01745_),
    .A2_N(_01751_),
    .B1(_01752_),
    .B2(_01746_),
    .X(_01773_));
 sky130_fd_sc_hd__o2111ai_2 _07863_ (.A1(_01585_),
    .A2(_01589_),
    .B1(_01591_),
    .C1(_01592_),
    .D1(_01588_),
    .Y(_01774_));
 sky130_fd_sc_hd__o21ai_1 _07864_ (.A1(_01587_),
    .A2(_01590_),
    .B1(_01593_),
    .Y(_01775_));
 sky130_fd_sc_hd__o21bai_1 _07865_ (.A1(_01587_),
    .A2(_01590_),
    .B1_N(_01593_),
    .Y(_01776_));
 sky130_fd_sc_hd__o211ai_1 _07866_ (.A1(_01585_),
    .A2(_01589_),
    .B1(_01588_),
    .C1(_01593_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand3_2 _07867_ (.A(_01773_),
    .B(_01774_),
    .C(_01775_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand3_2 _07868_ (.A(_01776_),
    .B(_01777_),
    .C(_01772_),
    .Y(_01779_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(net31),
    .B(net64),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _07870_ (.A(net31),
    .B(net34),
    .Y(_01781_));
 sky130_fd_sc_hd__nand4_2 _07871_ (.A(net32),
    .B(net31),
    .C(net64),
    .D(net34),
    .Y(_01783_));
 sky130_fd_sc_hd__a22oi_1 _07872_ (.A1(net32),
    .A2(net64),
    .B1(net34),
    .B2(net31),
    .Y(_01784_));
 sky130_fd_sc_hd__a22o_1 _07873_ (.A1(net32),
    .A2(net64),
    .B1(net34),
    .B2(net31),
    .X(_01785_));
 sky130_fd_sc_hd__and2_1 _07874_ (.A(net30),
    .B(net35),
    .X(_01786_));
 sky130_fd_sc_hd__nand2_1 _07875_ (.A(net30),
    .B(net35),
    .Y(_01787_));
 sky130_fd_sc_hd__o211ai_2 _07876_ (.A1(_01577_),
    .A2(_01780_),
    .B1(net30),
    .C1(_01785_),
    .Y(_01788_));
 sky130_fd_sc_hd__o211a_1 _07877_ (.A1(_01577_),
    .A2(_01780_),
    .B1(_01786_),
    .C1(_01785_),
    .X(_01789_));
 sky130_fd_sc_hd__o21ai_2 _07878_ (.A1(_01787_),
    .A2(_01784_),
    .B1(_01783_),
    .Y(_01790_));
 sky130_fd_sc_hd__o211ai_2 _07879_ (.A1(_00121_),
    .A2(_00407_),
    .B1(_01580_),
    .C1(_01581_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21oi_1 _07880_ (.A1(_01582_),
    .A2(_01791_),
    .B1(_01790_),
    .Y(_01792_));
 sky130_fd_sc_hd__a21o_1 _07881_ (.A1(_01582_),
    .A2(_01791_),
    .B1(_01790_),
    .X(_01794_));
 sky130_fd_sc_hd__and3_1 _07882_ (.A(_01582_),
    .B(_01790_),
    .C(_01791_),
    .X(_01795_));
 sky130_fd_sc_hd__nand3_1 _07883_ (.A(_01582_),
    .B(_01790_),
    .C(_01791_),
    .Y(_01796_));
 sky130_fd_sc_hd__o211ai_2 _07884_ (.A1(_01614_),
    .A2(_01615_),
    .B1(net28),
    .C1(net38),
    .Y(_01797_));
 sky130_fd_sc_hd__a211o_1 _07885_ (.A1(net28),
    .A2(net38),
    .B1(_01614_),
    .C1(_01615_),
    .X(_01798_));
 sky130_fd_sc_hd__nand2_1 _07886_ (.A(_01797_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21o_2 _07887_ (.A1(_01799_),
    .A2(_01794_),
    .B1(_01795_),
    .X(_01800_));
 sky130_fd_sc_hd__and3_1 _07888_ (.A(_01778_),
    .B(_01779_),
    .C(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__nand3_2 _07889_ (.A(_01778_),
    .B(_01779_),
    .C(_01800_),
    .Y(_01802_));
 sky130_fd_sc_hd__a21oi_2 _07890_ (.A1(_01778_),
    .A2(_01779_),
    .B1(_01800_),
    .Y(_01803_));
 sky130_fd_sc_hd__a21o_1 _07891_ (.A1(_01778_),
    .A2(_01779_),
    .B1(_01800_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _07892_ (.A(_01802_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__o21ai_1 _07893_ (.A1(_01801_),
    .A2(_01803_),
    .B1(_01769_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21boi_2 _07894_ (.A1(_01769_),
    .A2(_01806_),
    .B1_N(_01770_),
    .Y(_01808_));
 sky130_fd_sc_hd__nand4_2 _07895_ (.A(_01565_),
    .B(_01568_),
    .C(_01598_),
    .D(_01600_),
    .Y(_01809_));
 sky130_fd_sc_hd__o2bb2ai_4 _07896_ (.A1_N(_01565_),
    .A2_N(_01568_),
    .B1(_01597_),
    .B2(_01599_),
    .Y(_01810_));
 sky130_fd_sc_hd__a22oi_4 _07897_ (.A1(_01770_),
    .A2(_01807_),
    .B1(_01809_),
    .B2(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__o211a_1 _07898_ (.A1(_01567_),
    .A2(_01602_),
    .B1(_01808_),
    .C1(_01810_),
    .X(_01812_));
 sky130_fd_sc_hd__o211ai_2 _07899_ (.A1(_01567_),
    .A2(_01602_),
    .B1(_01808_),
    .C1(_01810_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21boi_1 _07900_ (.A1(_01778_),
    .A2(_01800_),
    .B1_N(_01779_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_01779_),
    .B(_01802_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand4_1 _07902_ (.A(_01643_),
    .B(_01644_),
    .C(_01657_),
    .D(_01658_),
    .Y(_01817_));
 sky130_fd_sc_hd__a22o_1 _07903_ (.A1(_01643_),
    .A2(_01644_),
    .B1(_01657_),
    .B2(_01658_),
    .X(_01818_));
 sky130_fd_sc_hd__o2bb2ai_1 _07904_ (.A1_N(_01643_),
    .A2_N(_01644_),
    .B1(_01655_),
    .B2(_01656_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand3_1 _07905_ (.A(_01659_),
    .B(_01644_),
    .C(_01643_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand3_1 _07906_ (.A(_01818_),
    .B(_01814_),
    .C(_01817_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand3_2 _07907_ (.A(_01816_),
    .B(_01819_),
    .C(_01820_),
    .Y(_01822_));
 sky130_fd_sc_hd__and4_1 _07908_ (.A(net28),
    .B(net29),
    .C(net37),
    .D(net36),
    .X(_01823_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(net27),
    .B(net38),
    .Y(_01824_));
 sky130_fd_sc_hd__a22oi_2 _07910_ (.A1(net28),
    .A2(net37),
    .B1(net36),
    .B2(net29),
    .Y(_01825_));
 sky130_fd_sc_hd__a22o_1 _07911_ (.A1(net28),
    .A2(net37),
    .B1(net36),
    .B2(net29),
    .X(_01827_));
 sky130_fd_sc_hd__and4b_1 _07912_ (.A_N(_01823_),
    .B(_01827_),
    .C(net27),
    .D(net38),
    .X(_01828_));
 sky130_fd_sc_hd__nand4b_1 _07913_ (.A_N(_01823_),
    .B(_01827_),
    .C(net27),
    .D(net38),
    .Y(_01829_));
 sky130_fd_sc_hd__o21bai_2 _07914_ (.A1(_01824_),
    .A2(_01825_),
    .B1_N(_01823_),
    .Y(_01830_));
 sky130_fd_sc_hd__a22oi_4 _07915_ (.A1(net23),
    .A2(net41),
    .B1(_01627_),
    .B2(_01629_),
    .Y(_01831_));
 sky130_fd_sc_hd__a22o_1 _07916_ (.A1(net23),
    .A2(net41),
    .B1(_01627_),
    .B2(_01629_),
    .X(_01832_));
 sky130_fd_sc_hd__o21bai_4 _07917_ (.A1(_01630_),
    .A2(_01831_),
    .B1_N(_01830_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _07918_ (.A(_01631_),
    .B(_01830_),
    .Y(_01834_));
 sky130_fd_sc_hd__nand3_1 _07919_ (.A(_01631_),
    .B(_01830_),
    .C(_01832_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _07920_ (.A(net23),
    .B(net39),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(net23),
    .B(net40),
    .Y(_01838_));
 sky130_fd_sc_hd__and4_1 _07922_ (.A(net26),
    .B(net23),
    .C(net39),
    .D(net40),
    .X(_01839_));
 sky130_fd_sc_hd__nand4_2 _07923_ (.A(net26),
    .B(net23),
    .C(net39),
    .D(net40),
    .Y(_01840_));
 sky130_fd_sc_hd__a22o_2 _07924_ (.A1(net26),
    .A2(net39),
    .B1(net40),
    .B2(net23),
    .X(_01841_));
 sky130_fd_sc_hd__o2111a_2 _07925_ (.A1(_01625_),
    .A2(_01836_),
    .B1(net12),
    .C1(net41),
    .D1(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__o2111ai_4 _07926_ (.A1(_01625_),
    .A2(_01836_),
    .B1(net12),
    .C1(net41),
    .D1(_01841_),
    .Y(_01843_));
 sky130_fd_sc_hd__a31o_1 _07927_ (.A1(_01841_),
    .A2(net41),
    .A3(net12),
    .B1(_01839_),
    .X(_01844_));
 sky130_fd_sc_hd__a31o_2 _07928_ (.A1(_01631_),
    .A2(_01830_),
    .A3(_01832_),
    .B1(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__o21ai_4 _07929_ (.A1(_01622_),
    .A2(_01633_),
    .B1(_01632_),
    .Y(_01846_));
 sky130_fd_sc_hd__a22oi_4 _07930_ (.A1(_01833_),
    .A2(_01845_),
    .B1(_01846_),
    .B2(_01636_),
    .Y(_01847_));
 sky130_fd_sc_hd__o2111a_1 _07931_ (.A1(_01622_),
    .A2(_01635_),
    .B1(_01833_),
    .C1(_01845_),
    .D1(_01846_),
    .X(_01849_));
 sky130_fd_sc_hd__o2111ai_4 _07932_ (.A1(_01622_),
    .A2(_01635_),
    .B1(_01833_),
    .C1(_01845_),
    .D1(_01846_),
    .Y(_01850_));
 sky130_fd_sc_hd__nand2_2 _07933_ (.A(net1),
    .B(net42),
    .Y(_01851_));
 sky130_fd_sc_hd__and4_1 _07934_ (.A(net12),
    .B(net1),
    .C(net43),
    .D(net42),
    .X(_01852_));
 sky130_fd_sc_hd__a22oi_2 _07935_ (.A1(net1),
    .A2(net45),
    .B1(_01646_),
    .B2(_01647_),
    .Y(_01853_));
 sky130_fd_sc_hd__or3b_2 _07936_ (.A(_01648_),
    .B(_01853_),
    .C_N(_01852_),
    .X(_01854_));
 sky130_fd_sc_hd__o32ai_2 _07937_ (.A1(_00022_),
    .A2(_00462_),
    .A3(_01851_),
    .B1(_01853_),
    .B2(_01648_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _07938_ (.A(_01854_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__o21ai_1 _07939_ (.A1(_01856_),
    .A2(_01847_),
    .B1(_01850_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21o_1 _07940_ (.A1(_01821_),
    .A2(_01822_),
    .B1(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__nand3_2 _07941_ (.A(_01821_),
    .B(_01822_),
    .C(_01857_),
    .Y(_01860_));
 sky130_fd_sc_hd__nand2_1 _07942_ (.A(_01858_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__a32oi_2 _07943_ (.A1(_01808_),
    .A2(_01809_),
    .A3(_01810_),
    .B1(_01858_),
    .B2(_01860_),
    .Y(_01862_));
 sky130_fd_sc_hd__o21ai_1 _07944_ (.A1(_01861_),
    .A2(_01811_),
    .B1(_01813_),
    .Y(_01863_));
 sky130_fd_sc_hd__nand3_1 _07945_ (.A(_01604_),
    .B(_01605_),
    .C(_01666_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21o_1 _07946_ (.A1(_01604_),
    .A2(_01605_),
    .B1(_01666_),
    .X(_01865_));
 sky130_fd_sc_hd__o2bb2ai_1 _07947_ (.A1_N(_01604_),
    .A2_N(_01605_),
    .B1(_01663_),
    .B2(_01665_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand4_1 _07948_ (.A(_01604_),
    .B(_01605_),
    .C(_01662_),
    .D(_01664_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand3_2 _07949_ (.A(_01866_),
    .B(_01867_),
    .C(_01863_),
    .Y(_01868_));
 sky130_fd_sc_hd__o211ai_2 _07950_ (.A1(_01811_),
    .A2(_01862_),
    .B1(_01864_),
    .C1(_01865_),
    .Y(_01869_));
 sky130_fd_sc_hd__o31a_1 _07951_ (.A1(_00033_),
    .A2(_00484_),
    .A3(_01654_),
    .B1(_01653_),
    .X(_01871_));
 sky130_fd_sc_hd__and2_1 _07952_ (.A(_01822_),
    .B(_01860_),
    .X(_01872_));
 sky130_fd_sc_hd__a21oi_1 _07953_ (.A1(_01822_),
    .A2(_01860_),
    .B1(_01871_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21o_2 _07954_ (.A1(_01822_),
    .A2(_01860_),
    .B1(_01871_),
    .X(_01874_));
 sky130_fd_sc_hd__o311a_1 _07955_ (.A1(_00033_),
    .A2(_00484_),
    .A3(_01654_),
    .B1(_01653_),
    .C1(_01872_),
    .X(_01875_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(_01871_),
    .B(_01872_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand4_2 _07957_ (.A(_01868_),
    .B(_01869_),
    .C(_01874_),
    .D(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__and2_2 _07958_ (.A(_01868_),
    .B(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__nand3_2 _07959_ (.A(_01671_),
    .B(_01674_),
    .C(_01681_),
    .Y(_01879_));
 sky130_fd_sc_hd__o21bai_2 _07960_ (.A1(_01670_),
    .A2(_01673_),
    .B1_N(_01681_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21ai_1 _07961_ (.A1(_01670_),
    .A2(_01673_),
    .B1(_01681_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand3_1 _07962_ (.A(_01671_),
    .B(_01674_),
    .C(_01680_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_1 _07963_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__a21oi_1 _07964_ (.A1(_01879_),
    .A2(_01880_),
    .B1(_01878_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand3b_2 _07965_ (.A_N(_01878_),
    .B(_01882_),
    .C(_01883_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand3_1 _07966_ (.A(_01880_),
    .B(_01878_),
    .C(_01879_),
    .Y(_01887_));
 sky130_fd_sc_hd__a31oi_4 _07967_ (.A1(_01880_),
    .A2(_01878_),
    .A3(_01879_),
    .B1(_01874_),
    .Y(_01888_));
 sky130_fd_sc_hd__a31o_1 _07968_ (.A1(_01880_),
    .A2(_01878_),
    .A3(_01879_),
    .B1(_01874_),
    .X(_01889_));
 sky130_fd_sc_hd__nand2_1 _07969_ (.A(_01690_),
    .B(_01692_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand3_1 _07970_ (.A(_01690_),
    .B(_01692_),
    .C(_01693_),
    .Y(_01891_));
 sky130_fd_sc_hd__o22ai_1 _07971_ (.A1(_01677_),
    .A2(_01679_),
    .B1(_01689_),
    .B2(_01691_),
    .Y(_01893_));
 sky130_fd_sc_hd__o211a_1 _07972_ (.A1(_01677_),
    .A2(_01679_),
    .B1(_01690_),
    .C1(_01692_),
    .X(_01894_));
 sky130_fd_sc_hd__o2bb2ai_1 _07973_ (.A1_N(_01693_),
    .A2_N(_01890_),
    .B1(_01888_),
    .B2(_01885_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _07974_ (.A(_01894_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__o2111ai_1 _07975_ (.A1(_01878_),
    .A2(_01884_),
    .B1(_01889_),
    .C1(_01891_),
    .D1(_01893_),
    .Y(_01897_));
 sky130_fd_sc_hd__o21a_2 _07976_ (.A1(_01894_),
    .A2(_01895_),
    .B1(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__o2bb2ai_2 _07977_ (.A1_N(_01868_),
    .A2_N(_01869_),
    .B1(_01873_),
    .B2(_01875_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand3b_1 _07978_ (.A_N(_01811_),
    .B(_01813_),
    .C(_01861_),
    .Y(_01900_));
 sky130_fd_sc_hd__o21bai_2 _07979_ (.A1(_01811_),
    .A2(_01812_),
    .B1_N(_01861_),
    .Y(_01901_));
 sky130_fd_sc_hd__o21ai_1 _07980_ (.A1(_01811_),
    .A2(_01812_),
    .B1(_01861_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand4b_1 _07981_ (.A_N(_01811_),
    .B(_01813_),
    .C(_01858_),
    .D(_01860_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_2 _07982_ (.A(net7),
    .B(net33),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_2 _07983_ (.A(net7),
    .B(net44),
    .Y(_01906_));
 sky130_fd_sc_hd__and4_1 _07984_ (.A(net7),
    .B(net8),
    .C(net44),
    .D(net33),
    .X(_01907_));
 sky130_fd_sc_hd__nand2_1 _07985_ (.A(net6),
    .B(net55),
    .Y(_01908_));
 sky130_fd_sc_hd__a22oi_4 _07986_ (.A1(net7),
    .A2(net44),
    .B1(net33),
    .B2(net8),
    .Y(_01909_));
 sky130_fd_sc_hd__a22o_1 _07987_ (.A1(net7),
    .A2(net44),
    .B1(net33),
    .B2(net8),
    .X(_01910_));
 sky130_fd_sc_hd__nand3_1 _07988_ (.A(_01906_),
    .B(net33),
    .C(net8),
    .Y(_01911_));
 sky130_fd_sc_hd__nand3_1 _07989_ (.A(_01703_),
    .B(net44),
    .C(net7),
    .Y(_01912_));
 sky130_fd_sc_hd__o2111ai_4 _07990_ (.A1(_01704_),
    .A2(_01905_),
    .B1(net6),
    .C1(net55),
    .D1(_01910_),
    .Y(_01913_));
 sky130_fd_sc_hd__o22ai_4 _07991_ (.A1(_01704_),
    .A2(_01905_),
    .B1(_01908_),
    .B2(_01909_),
    .Y(_01915_));
 sky130_fd_sc_hd__and3_1 _07992_ (.A(_01707_),
    .B(_01710_),
    .C(_01711_),
    .X(_01916_));
 sky130_fd_sc_hd__o211ai_4 _07993_ (.A1(_00176_),
    .A2(_00341_),
    .B1(_01710_),
    .C1(_01711_),
    .Y(_01917_));
 sky130_fd_sc_hd__o31a_1 _07994_ (.A1(_01707_),
    .A2(_01708_),
    .A3(_01706_),
    .B1(_01915_),
    .X(_01918_));
 sky130_fd_sc_hd__nand2_1 _07995_ (.A(_01712_),
    .B(_01915_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand3_2 _07996_ (.A(_01712_),
    .B(_01915_),
    .C(_01917_),
    .Y(_01920_));
 sky130_fd_sc_hd__a21oi_2 _07997_ (.A1(_01712_),
    .A2(_01917_),
    .B1(_01915_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21o_2 _07998_ (.A1(_01712_),
    .A2(_01917_),
    .B1(_01915_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(net4),
    .B(net60),
    .Y(_01923_));
 sky130_fd_sc_hd__nand4_4 _08000_ (.A(net5),
    .B(net6),
    .C(net58),
    .D(net59),
    .Y(_01924_));
 sky130_fd_sc_hd__o22a_1 _08001_ (.A1(_00187_),
    .A2(_00330_),
    .B1(_00363_),
    .B2(_00154_),
    .X(_01926_));
 sky130_fd_sc_hd__a22o_2 _08002_ (.A1(net6),
    .A2(net58),
    .B1(net59),
    .B2(net5),
    .X(_01927_));
 sky130_fd_sc_hd__o211ai_2 _08003_ (.A1(_00165_),
    .A2(_00352_),
    .B1(_01924_),
    .C1(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__a21o_1 _08004_ (.A1(_01924_),
    .A2(_01927_),
    .B1(_01923_),
    .X(_01929_));
 sky130_fd_sc_hd__o2bb2a_1 _08005_ (.A1_N(_01924_),
    .A2_N(_01927_),
    .B1(_00165_),
    .B2(_00352_),
    .X(_01930_));
 sky130_fd_sc_hd__a22o_1 _08006_ (.A1(net4),
    .A2(net60),
    .B1(_01924_),
    .B2(_01927_),
    .X(_01931_));
 sky130_fd_sc_hd__and4_1 _08007_ (.A(_01927_),
    .B(net60),
    .C(net4),
    .D(_01924_),
    .X(_01932_));
 sky130_fd_sc_hd__nand4_2 _08008_ (.A(_01927_),
    .B(net60),
    .C(net4),
    .D(_01924_),
    .Y(_01933_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_01931_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__a221oi_4 _08010_ (.A1(_01928_),
    .A2(_01929_),
    .B1(_01918_),
    .B2(_01917_),
    .C1(_01921_),
    .Y(_01935_));
 sky130_fd_sc_hd__o2111ai_4 _08011_ (.A1(_01919_),
    .A2(_01916_),
    .B1(_01931_),
    .C1(_01922_),
    .D1(_01933_),
    .Y(_01937_));
 sky130_fd_sc_hd__o22a_2 _08012_ (.A1(_01916_),
    .A2(_01919_),
    .B1(_01921_),
    .B2(_01934_),
    .X(_01938_));
 sky130_fd_sc_hd__o21ai_1 _08013_ (.A1(_01921_),
    .A2(_01934_),
    .B1(_01920_),
    .Y(_01939_));
 sky130_fd_sc_hd__o211ai_4 _08014_ (.A1(_01724_),
    .A2(_01725_),
    .B1(_01729_),
    .C1(_01717_),
    .Y(_01940_));
 sky130_fd_sc_hd__o2bb2ai_4 _08015_ (.A1_N(_01722_),
    .A2_N(_01723_),
    .B1(_01728_),
    .B2(_01715_),
    .Y(_01941_));
 sky130_fd_sc_hd__o22ai_1 _08016_ (.A1(_01724_),
    .A2(_01725_),
    .B1(_01728_),
    .B2(_01715_),
    .Y(_01942_));
 sky130_fd_sc_hd__a21oi_4 _08017_ (.A1(_01940_),
    .A2(_01941_),
    .B1(_01938_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand3_2 _08018_ (.A(_01732_),
    .B(_01939_),
    .C(_01942_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand3_4 _08019_ (.A(_01938_),
    .B(_01940_),
    .C(_01941_),
    .Y(_01945_));
 sky130_fd_sc_hd__nand2_2 _08020_ (.A(net2),
    .B(net61),
    .Y(_01946_));
 sky130_fd_sc_hd__and4_1 _08021_ (.A(net3),
    .B(net2),
    .C(net62),
    .D(net61),
    .X(_01948_));
 sky130_fd_sc_hd__nand4_1 _08022_ (.A(net3),
    .B(net2),
    .C(net62),
    .D(net61),
    .Y(_01949_));
 sky130_fd_sc_hd__a22o_2 _08023_ (.A1(net2),
    .A2(net62),
    .B1(net61),
    .B2(net3),
    .X(_01950_));
 sky130_fd_sc_hd__and4_1 _08024_ (.A(_01950_),
    .B(net63),
    .C(net32),
    .D(_01949_),
    .X(_01951_));
 sky130_fd_sc_hd__o2111ai_4 _08025_ (.A1(_01737_),
    .A2(_01946_),
    .B1(net32),
    .C1(net63),
    .D1(_01950_),
    .Y(_01952_));
 sky130_fd_sc_hd__a31o_1 _08026_ (.A1(_01950_),
    .A2(net63),
    .A3(net32),
    .B1(_01948_),
    .X(_01953_));
 sky130_fd_sc_hd__o211ai_2 _08027_ (.A1(_00143_),
    .A2(_00396_),
    .B1(_01741_),
    .C1(_01742_),
    .Y(_01954_));
 sky130_fd_sc_hd__o21a_1 _08028_ (.A1(_00165_),
    .A2(_00352_),
    .B1(_01924_),
    .X(_01955_));
 sky130_fd_sc_hd__o21ai_1 _08029_ (.A1(_00165_),
    .A2(_00352_),
    .B1(_01924_),
    .Y(_01956_));
 sky130_fd_sc_hd__nand4_2 _08030_ (.A(_01743_),
    .B(_01927_),
    .C(_01954_),
    .D(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__o2bb2ai_2 _08031_ (.A1_N(_01743_),
    .A2_N(_01954_),
    .B1(_01955_),
    .B2(_01926_),
    .Y(_01959_));
 sky130_fd_sc_hd__o211a_1 _08032_ (.A1(_01948_),
    .A2(_01951_),
    .B1(_01957_),
    .C1(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__a21oi_2 _08033_ (.A1(_01957_),
    .A2(_01959_),
    .B1(_01953_),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_2 _08034_ (.A(_01960_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_2 _08035_ (.A(_01945_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_2 _08036_ (.A1(_01945_),
    .A2(_01962_),
    .B1(_01943_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21o_1 _08037_ (.A1(_01945_),
    .A2(_01962_),
    .B1(_01943_),
    .X(_01965_));
 sky130_fd_sc_hd__a221o_1 _08038_ (.A1(_01717_),
    .A2(_01732_),
    .B1(_01755_),
    .B2(_01757_),
    .C1(_01702_),
    .X(_01966_));
 sky130_fd_sc_hd__o211ai_1 _08039_ (.A1(_01728_),
    .A2(_01731_),
    .B1(_01759_),
    .C1(_01702_),
    .Y(_01967_));
 sky130_fd_sc_hd__o211ai_2 _08040_ (.A1(_01733_),
    .A2(_01702_),
    .B1(_01967_),
    .C1(_01762_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _08041_ (.A(_01735_),
    .B(_01736_),
    .Y(_01970_));
 sky130_fd_sc_hd__o21ai_1 _08042_ (.A1(_01702_),
    .A2(_01733_),
    .B1(_01761_),
    .Y(_01971_));
 sky130_fd_sc_hd__a21o_1 _08043_ (.A1(_01735_),
    .A2(_01736_),
    .B1(_01758_),
    .X(_01972_));
 sky130_fd_sc_hd__and3_1 _08044_ (.A(_01968_),
    .B(_01964_),
    .C(_01966_),
    .X(_01973_));
 sky130_fd_sc_hd__nand3_2 _08045_ (.A(_01968_),
    .B(_01964_),
    .C(_01966_),
    .Y(_01974_));
 sky130_fd_sc_hd__a22oi_1 _08046_ (.A1(_01944_),
    .A2(_01963_),
    .B1(_01970_),
    .B2(_01759_),
    .Y(_01975_));
 sky130_fd_sc_hd__o211a_1 _08047_ (.A1(_01734_),
    .A2(_01762_),
    .B1(_01965_),
    .C1(_01972_),
    .X(_01976_));
 sky130_fd_sc_hd__o211ai_4 _08048_ (.A1(_01734_),
    .A2(_01762_),
    .B1(_01965_),
    .C1(_01972_),
    .Y(_01977_));
 sky130_fd_sc_hd__a21boi_4 _08049_ (.A1(_01953_),
    .A2(_01959_),
    .B1_N(_01957_),
    .Y(_01978_));
 sky130_fd_sc_hd__o21ai_2 _08050_ (.A1(_01792_),
    .A2(_01795_),
    .B1(_01799_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand4_2 _08051_ (.A(_01794_),
    .B(_01796_),
    .C(_01797_),
    .D(_01798_),
    .Y(_01981_));
 sky130_fd_sc_hd__nand3_1 _08052_ (.A(_01799_),
    .B(_01796_),
    .C(_01794_),
    .Y(_01982_));
 sky130_fd_sc_hd__a21o_1 _08053_ (.A1(_01794_),
    .A2(_01796_),
    .B1(_01799_),
    .X(_01983_));
 sky130_fd_sc_hd__a21oi_1 _08054_ (.A1(_01979_),
    .A2(_01981_),
    .B1(_01978_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand3b_4 _08055_ (.A_N(_01978_),
    .B(_01982_),
    .C(_01983_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand3_4 _08056_ (.A(_01978_),
    .B(_01979_),
    .C(_01981_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(net30),
    .B(net64),
    .Y(_01987_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(net30),
    .B(net34),
    .Y(_01988_));
 sky130_fd_sc_hd__and2_1 _08059_ (.A(net29),
    .B(net35),
    .X(_01989_));
 sky130_fd_sc_hd__a22o_1 _08060_ (.A1(net31),
    .A2(net64),
    .B1(net34),
    .B2(net30),
    .X(_01990_));
 sky130_fd_sc_hd__nand3_1 _08061_ (.A(_01988_),
    .B(net64),
    .C(net31),
    .Y(_01992_));
 sky130_fd_sc_hd__nand3_1 _08062_ (.A(_01780_),
    .B(net34),
    .C(net30),
    .Y(_01993_));
 sky130_fd_sc_hd__o2111ai_4 _08063_ (.A1(_01781_),
    .A2(_01987_),
    .B1(net29),
    .C1(net35),
    .D1(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__o2bb2ai_2 _08064_ (.A1_N(_01989_),
    .A2_N(_01990_),
    .B1(_01781_),
    .B2(_01987_),
    .Y(_01995_));
 sky130_fd_sc_hd__a21oi_1 _08065_ (.A1(_01783_),
    .A2(_01785_),
    .B1(_01786_),
    .Y(_01996_));
 sky130_fd_sc_hd__a22o_1 _08066_ (.A1(net30),
    .A2(net35),
    .B1(_01783_),
    .B2(_01785_),
    .X(_01997_));
 sky130_fd_sc_hd__o211ai_4 _08067_ (.A1(_00407_),
    .A2(_01788_),
    .B1(_01995_),
    .C1(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o221a_2 _08068_ (.A1(_01780_),
    .A2(_01988_),
    .B1(_01996_),
    .B2(_01789_),
    .C1(_01994_),
    .X(_01999_));
 sky130_fd_sc_hd__o21bai_2 _08069_ (.A1(_01789_),
    .A2(_01996_),
    .B1_N(_01995_),
    .Y(_02000_));
 sky130_fd_sc_hd__o2bb2a_1 _08070_ (.A1_N(net27),
    .A2_N(net38),
    .B1(_01823_),
    .B2(_01825_),
    .X(_02001_));
 sky130_fd_sc_hd__o21ai_1 _08071_ (.A1(_01823_),
    .A2(_01825_),
    .B1(_01824_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_2 _08072_ (.A(_01829_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__o21a_1 _08073_ (.A1(_01828_),
    .A2(_02001_),
    .B1(_01998_),
    .X(_02005_));
 sky130_fd_sc_hd__a21oi_2 _08074_ (.A1(_01998_),
    .A2(_02004_),
    .B1(_01999_),
    .Y(_02006_));
 sky130_fd_sc_hd__o211a_1 _08075_ (.A1(_01999_),
    .A2(_02005_),
    .B1(_01985_),
    .C1(_01986_),
    .X(_02007_));
 sky130_fd_sc_hd__a221oi_4 _08076_ (.A1(_01985_),
    .A2(_01986_),
    .B1(_01998_),
    .B2(_02004_),
    .C1(_01999_),
    .Y(_02008_));
 sky130_fd_sc_hd__o2bb2a_1 _08077_ (.A1_N(_01985_),
    .A2_N(_01986_),
    .B1(_01999_),
    .B2(_02005_),
    .X(_02009_));
 sky130_fd_sc_hd__o2bb2ai_2 _08078_ (.A1_N(_01985_),
    .A2_N(_01986_),
    .B1(_01999_),
    .B2(_02005_),
    .Y(_02010_));
 sky130_fd_sc_hd__and3_1 _08079_ (.A(_01985_),
    .B(_01986_),
    .C(_02006_),
    .X(_02011_));
 sky130_fd_sc_hd__nand3_2 _08080_ (.A(_01985_),
    .B(_01986_),
    .C(_02006_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_02010_),
    .B(_02012_),
    .Y(_02014_));
 sky130_fd_sc_hd__a22oi_2 _08082_ (.A1(_02010_),
    .A2(_02012_),
    .B1(_01975_),
    .B2(_01971_),
    .Y(_02015_));
 sky130_fd_sc_hd__a31oi_2 _08083_ (.A1(_01966_),
    .A2(_01968_),
    .A3(_01964_),
    .B1(_02014_),
    .Y(_02016_));
 sky130_fd_sc_hd__a21o_1 _08084_ (.A1(_01769_),
    .A2(_01770_),
    .B1(_01806_),
    .X(_02017_));
 sky130_fd_sc_hd__o211ai_1 _08085_ (.A1(_01801_),
    .A2(_01803_),
    .B1(_01769_),
    .C1(_01770_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand4_4 _08086_ (.A(_01769_),
    .B(_01770_),
    .C(_01802_),
    .D(_01805_),
    .Y(_02019_));
 sky130_fd_sc_hd__o2bb2ai_2 _08087_ (.A1_N(_01769_),
    .A2_N(_01770_),
    .B1(_01801_),
    .B2(_01803_),
    .Y(_02020_));
 sky130_fd_sc_hd__a2bb2oi_2 _08088_ (.A1_N(_01973_),
    .A2_N(_02015_),
    .B1(_02019_),
    .B2(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__o211ai_2 _08089_ (.A1(_01973_),
    .A2(_02015_),
    .B1(_02017_),
    .C1(_02018_),
    .Y(_02022_));
 sky130_fd_sc_hd__o211a_1 _08090_ (.A1(_01976_),
    .A2(_02016_),
    .B1(_02019_),
    .C1(_02020_),
    .X(_02023_));
 sky130_fd_sc_hd__o211ai_4 _08091_ (.A1(_01976_),
    .A2(_02016_),
    .B1(_02019_),
    .C1(_02020_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(net27),
    .B(net37),
    .Y(_02026_));
 sky130_fd_sc_hd__a22oi_4 _08093_ (.A1(net27),
    .A2(net37),
    .B1(net36),
    .B2(net28),
    .Y(_02027_));
 sky130_fd_sc_hd__a22o_1 _08094_ (.A1(net27),
    .A2(net37),
    .B1(net36),
    .B2(net28),
    .X(_02028_));
 sky130_fd_sc_hd__nand4_4 _08095_ (.A(net28),
    .B(net27),
    .C(net37),
    .D(net36),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _08096_ (.A(net26),
    .B(net38),
    .Y(_02030_));
 sky130_fd_sc_hd__and2_1 _08097_ (.A(_02029_),
    .B(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__o21ai_1 _08098_ (.A1(_02030_),
    .A2(_02027_),
    .B1(_02029_),
    .Y(_02032_));
 sky130_fd_sc_hd__a2bb2oi_2 _08099_ (.A1_N(_00022_),
    .A2_N(_00451_),
    .B1(_01840_),
    .B2(_01841_),
    .Y(_02033_));
 sky130_fd_sc_hd__a22o_1 _08100_ (.A1(net12),
    .A2(net41),
    .B1(_01840_),
    .B2(_01841_),
    .X(_02034_));
 sky130_fd_sc_hd__nand2_1 _08101_ (.A(_02032_),
    .B(_01843_),
    .Y(_02036_));
 sky130_fd_sc_hd__and3_2 _08102_ (.A(_01843_),
    .B(_02034_),
    .C(_02032_),
    .X(_02037_));
 sky130_fd_sc_hd__nand3_1 _08103_ (.A(_01843_),
    .B(_02034_),
    .C(_02032_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _08104_ (.A(net12),
    .B(net39),
    .Y(_02039_));
 sky130_fd_sc_hd__and4_1 _08105_ (.A(net12),
    .B(net23),
    .C(net39),
    .D(net40),
    .X(_02040_));
 sky130_fd_sc_hd__a22oi_1 _08106_ (.A1(net23),
    .A2(net39),
    .B1(net40),
    .B2(net12),
    .Y(_02041_));
 sky130_fd_sc_hd__a22o_1 _08107_ (.A1(net23),
    .A2(net39),
    .B1(net40),
    .B2(net12),
    .X(_02042_));
 sky130_fd_sc_hd__o2111a_1 _08108_ (.A1(_01838_),
    .A2(_02039_),
    .B1(net1),
    .C1(net41),
    .D1(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__o2111ai_2 _08109_ (.A1(_01838_),
    .A2(_02039_),
    .B1(net1),
    .C1(net41),
    .D1(_02042_),
    .Y(_02044_));
 sky130_fd_sc_hd__a31o_1 _08110_ (.A1(_02042_),
    .A2(net41),
    .A3(net1),
    .B1(_02040_),
    .X(_02045_));
 sky130_fd_sc_hd__o22ai_4 _08111_ (.A1(_02027_),
    .A2(_02031_),
    .B1(_02033_),
    .B2(_01842_),
    .Y(_02047_));
 sky130_fd_sc_hd__o21ai_1 _08112_ (.A1(_02040_),
    .A2(_02043_),
    .B1(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__o221a_2 _08113_ (.A1(_02040_),
    .A2(_02043_),
    .B1(_02033_),
    .B2(_02036_),
    .C1(_02047_),
    .X(_02049_));
 sky130_fd_sc_hd__o2bb2a_1 _08114_ (.A1_N(_02045_),
    .A2_N(_02047_),
    .B1(_02033_),
    .B2(_02036_),
    .X(_02050_));
 sky130_fd_sc_hd__a22o_1 _08115_ (.A1(_01833_),
    .A2(_01835_),
    .B1(_01840_),
    .B2(_01843_),
    .X(_02051_));
 sky130_fd_sc_hd__o2111ai_1 _08116_ (.A1(_01625_),
    .A2(_01836_),
    .B1(_01843_),
    .C1(_01833_),
    .D1(_01835_),
    .Y(_02052_));
 sky130_fd_sc_hd__o221ai_4 _08117_ (.A1(_01839_),
    .A2(_01842_),
    .B1(_01831_),
    .B2(_01834_),
    .C1(_01833_),
    .Y(_02053_));
 sky130_fd_sc_hd__a21o_1 _08118_ (.A1(_01833_),
    .A2(_01835_),
    .B1(_01844_),
    .X(_02054_));
 sky130_fd_sc_hd__o211ai_4 _08119_ (.A1(_02037_),
    .A2(_02049_),
    .B1(_02053_),
    .C1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand3_2 _08120_ (.A(_02051_),
    .B(_02052_),
    .C(_02050_),
    .Y(_02056_));
 sky130_fd_sc_hd__o22a_1 _08121_ (.A1(_00033_),
    .A2(_00462_),
    .B1(_00473_),
    .B2(_00022_),
    .X(_02058_));
 sky130_fd_sc_hd__o211a_1 _08122_ (.A1(_00033_),
    .A2(_00462_),
    .B1(net42),
    .C1(net12),
    .X(_02059_));
 sky130_fd_sc_hd__o211a_1 _08123_ (.A1(_00022_),
    .A2(_00473_),
    .B1(net43),
    .C1(net1),
    .X(_02060_));
 sky130_fd_sc_hd__o21ai_1 _08124_ (.A1(_01852_),
    .A2(_02058_),
    .B1(_02055_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _08125_ (.A(_02056_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand3b_1 _08126_ (.A_N(_01847_),
    .B(_01850_),
    .C(_01856_),
    .Y(_02063_));
 sky130_fd_sc_hd__o21bai_1 _08127_ (.A1(_01847_),
    .A2(_01849_),
    .B1_N(_01856_),
    .Y(_02064_));
 sky130_fd_sc_hd__o21ai_1 _08128_ (.A1(_01847_),
    .A2(_01849_),
    .B1(_01856_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand4b_1 _08129_ (.A_N(_01847_),
    .B(_01850_),
    .C(_01854_),
    .D(_01855_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21o_1 _08130_ (.A1(_01986_),
    .A2(_02006_),
    .B1(_01984_),
    .X(_02067_));
 sky130_fd_sc_hd__a21oi_1 _08131_ (.A1(_01986_),
    .A2(_02006_),
    .B1(_01984_),
    .Y(_02069_));
 sky130_fd_sc_hd__and3_1 _08132_ (.A(_02063_),
    .B(_02064_),
    .C(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__nand3_1 _08133_ (.A(_02063_),
    .B(_02064_),
    .C(_02069_),
    .Y(_02071_));
 sky130_fd_sc_hd__nand3_1 _08134_ (.A(_02065_),
    .B(_02066_),
    .C(_02067_),
    .Y(_02072_));
 sky130_fd_sc_hd__a31o_1 _08135_ (.A1(_02065_),
    .A2(_02066_),
    .A3(_02067_),
    .B1(_02062_),
    .X(_02073_));
 sky130_fd_sc_hd__a22o_1 _08136_ (.A1(_02056_),
    .A2(_02061_),
    .B1(_02071_),
    .B2(_02072_),
    .X(_02074_));
 sky130_fd_sc_hd__o21ai_4 _08137_ (.A1(_02070_),
    .A2(_02073_),
    .B1(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__o21ai_1 _08138_ (.A1(_02021_),
    .A2(_02075_),
    .B1(_02025_),
    .Y(_02076_));
 sky130_fd_sc_hd__o2111ai_4 _08139_ (.A1(_02021_),
    .A2(_02075_),
    .B1(_02025_),
    .C1(_01900_),
    .D1(_01901_),
    .Y(_02077_));
 sky130_fd_sc_hd__inv_2 _08140_ (.A(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_1 _08141_ (.A(_01902_),
    .B(_01904_),
    .C(_02076_),
    .Y(_02080_));
 sky130_fd_sc_hd__o21a_1 _08142_ (.A1(_02070_),
    .A2(_02073_),
    .B1(_02072_),
    .X(_02081_));
 sky130_fd_sc_hd__nor2_1 _08143_ (.A(_01854_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__xnor2_1 _08144_ (.A(_01854_),
    .B(_02081_),
    .Y(_02083_));
 sky130_fd_sc_hd__and2_1 _08145_ (.A(_02080_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__nand2_1 _08146_ (.A(_02080_),
    .B(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand4_4 _08147_ (.A(_01877_),
    .B(_01899_),
    .C(_02077_),
    .D(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__o2bb2ai_1 _08148_ (.A1_N(_01877_),
    .A2_N(_01899_),
    .B1(_02078_),
    .B2(_02084_),
    .Y(_02087_));
 sky130_fd_sc_hd__nand3_2 _08149_ (.A(_02087_),
    .B(_02082_),
    .C(_02086_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_2 _08150_ (.A(_02086_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_01886_),
    .B(_01887_),
    .Y(_02091_));
 sky130_fd_sc_hd__a22oi_4 _08152_ (.A1(_01886_),
    .A2(_01888_),
    .B1(_02091_),
    .B2(_01874_),
    .Y(_02092_));
 sky130_fd_sc_hd__o2bb2ai_1 _08153_ (.A1_N(_01874_),
    .A2_N(_02091_),
    .B1(_01889_),
    .B2(_01885_),
    .Y(_02093_));
 sky130_fd_sc_hd__nand3_1 _08154_ (.A(_02086_),
    .B(_02088_),
    .C(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_2 _08155_ (.A(net4),
    .B(net44),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_2 _08156_ (.A(net3),
    .B(net33),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_2 _08157_ (.A(net4),
    .B(net33),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _08158_ (.A(net3),
    .B(net44),
    .Y(_02098_));
 sky130_fd_sc_hd__and2_1 _08159_ (.A(net2),
    .B(net55),
    .X(_02099_));
 sky130_fd_sc_hd__nand2_1 _08160_ (.A(net2),
    .B(net55),
    .Y(_02100_));
 sky130_fd_sc_hd__a22oi_2 _08161_ (.A1(net3),
    .A2(net44),
    .B1(net33),
    .B2(net4),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _08162_ (.A(_02097_),
    .B(_02098_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand3_1 _08163_ (.A(_02098_),
    .B(net33),
    .C(net4),
    .Y(_02104_));
 sky130_fd_sc_hd__nand3_1 _08164_ (.A(_02097_),
    .B(net44),
    .C(net3),
    .Y(_02105_));
 sky130_fd_sc_hd__o211ai_4 _08165_ (.A1(_02095_),
    .A2(_02096_),
    .B1(_02099_),
    .C1(_02103_),
    .Y(_02106_));
 sky130_fd_sc_hd__o22ai_4 _08166_ (.A1(_02095_),
    .A2(_02096_),
    .B1(_02100_),
    .B2(_02102_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(net5),
    .B(net44),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_2 _08168_ (.A(net5),
    .B(net33),
    .Y(_02109_));
 sky130_fd_sc_hd__nand4_4 _08169_ (.A(net5),
    .B(net4),
    .C(net44),
    .D(net33),
    .Y(_02110_));
 sky130_fd_sc_hd__a22oi_1 _08170_ (.A1(net4),
    .A2(net44),
    .B1(net33),
    .B2(net5),
    .Y(_02111_));
 sky130_fd_sc_hd__a22o_2 _08171_ (.A1(net4),
    .A2(net44),
    .B1(net33),
    .B2(net5),
    .X(_02113_));
 sky130_fd_sc_hd__and2_1 _08172_ (.A(net3),
    .B(net55),
    .X(_02114_));
 sky130_fd_sc_hd__nand2_1 _08173_ (.A(net3),
    .B(net55),
    .Y(_02115_));
 sky130_fd_sc_hd__o211a_1 _08174_ (.A1(_02097_),
    .A2(_02108_),
    .B1(_02114_),
    .C1(_02113_),
    .X(_02116_));
 sky130_fd_sc_hd__o2111ai_4 _08175_ (.A1(_02097_),
    .A2(_02108_),
    .B1(net3),
    .C1(net55),
    .D1(_02113_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21oi_4 _08176_ (.A1(_02110_),
    .A2(_02113_),
    .B1(_02114_),
    .Y(_02118_));
 sky130_fd_sc_hd__o2bb2ai_1 _08177_ (.A1_N(_02110_),
    .A2_N(_02113_),
    .B1(_00132_),
    .B2(_00341_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_2 _08178_ (.A(_02107_),
    .B(_02117_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand3_1 _08179_ (.A(_02107_),
    .B(_02117_),
    .C(_02119_),
    .Y(_02121_));
 sky130_fd_sc_hd__a21oi_1 _08180_ (.A1(_02117_),
    .A2(_02119_),
    .B1(_02107_),
    .Y(_02122_));
 sky130_fd_sc_hd__o21bai_4 _08181_ (.A1(_02116_),
    .A2(_02118_),
    .B1_N(_02107_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_1 _08182_ (.A(net31),
    .B(net60),
    .Y(_02125_));
 sky130_fd_sc_hd__a22oi_4 _08183_ (.A1(net2),
    .A2(net58),
    .B1(net59),
    .B2(net32),
    .Y(_02126_));
 sky130_fd_sc_hd__and4_1 _08184_ (.A(net32),
    .B(net2),
    .C(net58),
    .D(net59),
    .X(_02127_));
 sky130_fd_sc_hd__nand4_1 _08185_ (.A(net32),
    .B(net2),
    .C(net58),
    .D(net59),
    .Y(_02128_));
 sky130_fd_sc_hd__a211oi_2 _08186_ (.A1(net31),
    .A2(net60),
    .B1(_02126_),
    .C1(_02127_),
    .Y(_02129_));
 sky130_fd_sc_hd__o211a_1 _08187_ (.A1(_02126_),
    .A2(_02127_),
    .B1(net31),
    .C1(net60),
    .X(_02130_));
 sky130_fd_sc_hd__o22a_1 _08188_ (.A1(_00121_),
    .A2(_00352_),
    .B1(_02126_),
    .B2(_02127_),
    .X(_02131_));
 sky130_fd_sc_hd__and4b_1 _08189_ (.A_N(_02126_),
    .B(_02128_),
    .C(net31),
    .D(net60),
    .X(_02132_));
 sky130_fd_sc_hd__nor2_1 _08190_ (.A(_02129_),
    .B(_02130_),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _08191_ (.A(_02131_),
    .B(_02132_),
    .Y(_02135_));
 sky130_fd_sc_hd__o221a_1 _08192_ (.A1(_02118_),
    .A2(_02120_),
    .B1(_02129_),
    .B2(_02130_),
    .C1(_02124_),
    .X(_02136_));
 sky130_fd_sc_hd__o221ai_4 _08193_ (.A1(_02118_),
    .A2(_02120_),
    .B1(_02129_),
    .B2(_02130_),
    .C1(_02124_),
    .Y(_02137_));
 sky130_fd_sc_hd__o22ai_4 _08194_ (.A1(_02118_),
    .A2(_02120_),
    .B1(_02122_),
    .B2(_02133_),
    .Y(_02138_));
 sky130_fd_sc_hd__o21ai_2 _08195_ (.A1(_02115_),
    .A2(_02111_),
    .B1(_02110_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _08196_ (.A(net4),
    .B(net55),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_2 _08197_ (.A(net6),
    .B(net44),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_2 _08198_ (.A(net6),
    .B(net33),
    .Y(_02142_));
 sky130_fd_sc_hd__a22oi_2 _08199_ (.A1(net5),
    .A2(net44),
    .B1(net33),
    .B2(net6),
    .Y(_02143_));
 sky130_fd_sc_hd__a22o_1 _08200_ (.A1(net5),
    .A2(net44),
    .B1(net33),
    .B2(net6),
    .X(_02144_));
 sky130_fd_sc_hd__nand3_1 _08201_ (.A(_02108_),
    .B(net33),
    .C(net6),
    .Y(_02146_));
 sky130_fd_sc_hd__nand3_1 _08202_ (.A(_02142_),
    .B(net44),
    .C(net5),
    .Y(_02147_));
 sky130_fd_sc_hd__o2111ai_4 _08203_ (.A1(_02109_),
    .A2(_02141_),
    .B1(net4),
    .C1(net55),
    .D1(_02144_),
    .Y(_02148_));
 sky130_fd_sc_hd__and3_2 _08204_ (.A(_02140_),
    .B(_02146_),
    .C(_02147_),
    .X(_02149_));
 sky130_fd_sc_hd__o211ai_1 _08205_ (.A1(_00165_),
    .A2(_00341_),
    .B1(_02146_),
    .C1(_02147_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_2 _08206_ (.A(_02139_),
    .B(_02148_),
    .Y(_02151_));
 sky130_fd_sc_hd__nand3_1 _08207_ (.A(_02139_),
    .B(_02148_),
    .C(_02150_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21o_2 _08208_ (.A1(_02148_),
    .A2(_02150_),
    .B1(_02139_),
    .X(_02153_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(net32),
    .B(net60),
    .Y(_02154_));
 sky130_fd_sc_hd__a22oi_2 _08210_ (.A1(net3),
    .A2(net58),
    .B1(net59),
    .B2(net2),
    .Y(_02155_));
 sky130_fd_sc_hd__a22o_1 _08211_ (.A1(net3),
    .A2(net58),
    .B1(net59),
    .B2(net2),
    .X(_02157_));
 sky130_fd_sc_hd__nand4_2 _08212_ (.A(net3),
    .B(net2),
    .C(net58),
    .D(net59),
    .Y(_02158_));
 sky130_fd_sc_hd__a22oi_2 _08213_ (.A1(net32),
    .A2(net60),
    .B1(_02157_),
    .B2(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor3b_1 _08214_ (.A(_02154_),
    .B(_02155_),
    .C_N(_02158_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_2 _08215_ (.A(_02159_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__o211ai_4 _08216_ (.A1(_02151_),
    .A2(_02149_),
    .B1(_02161_),
    .C1(_02153_),
    .Y(_02162_));
 sky130_fd_sc_hd__inv_2 _08217_ (.A(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__o2bb2ai_2 _08218_ (.A1_N(_02152_),
    .A2_N(_02153_),
    .B1(_02159_),
    .B2(_02160_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_2 _08219_ (.A1(_02162_),
    .A2(_02164_),
    .B1(_02138_),
    .Y(_02165_));
 sky130_fd_sc_hd__a21o_2 _08220_ (.A1(_02162_),
    .A2(_02164_),
    .B1(_02138_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_2 _08221_ (.A(_02138_),
    .B(_02164_),
    .Y(_02168_));
 sky130_fd_sc_hd__and3_1 _08222_ (.A(_02138_),
    .B(_02162_),
    .C(_02164_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_4 _08223_ (.A(net30),
    .B(net62),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_2 _08224_ (.A(net29),
    .B(net61),
    .Y(_02171_));
 sky130_fd_sc_hd__nand2_1 _08225_ (.A(net30),
    .B(net61),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _08226_ (.A(net29),
    .B(net62),
    .Y(_02173_));
 sky130_fd_sc_hd__nand4_1 _08227_ (.A(net30),
    .B(net29),
    .C(net62),
    .D(net61),
    .Y(_02174_));
 sky130_fd_sc_hd__a22o_2 _08228_ (.A1(net29),
    .A2(net62),
    .B1(net61),
    .B2(net30),
    .X(_02175_));
 sky130_fd_sc_hd__o211ai_4 _08229_ (.A1(_02170_),
    .A2(_02171_),
    .B1(net63),
    .C1(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__o2111ai_4 _08230_ (.A1(_02170_),
    .A2(_02171_),
    .B1(net28),
    .C1(net63),
    .D1(_02175_),
    .Y(_02177_));
 sky130_fd_sc_hd__o31a_2 _08231_ (.A1(_00088_),
    .A2(_00374_),
    .A3(_02171_),
    .B1(_02177_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _08232_ (.A(net31),
    .B(net62),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_4 _08233_ (.A(net31),
    .B(net61),
    .Y(_02181_));
 sky130_fd_sc_hd__a22o_1 _08234_ (.A1(net30),
    .A2(net62),
    .B1(net61),
    .B2(net31),
    .X(_02182_));
 sky130_fd_sc_hd__nand3_1 _08235_ (.A(_02170_),
    .B(net61),
    .C(net31),
    .Y(_02183_));
 sky130_fd_sc_hd__nand3_1 _08236_ (.A(_02181_),
    .B(net62),
    .C(net30),
    .Y(_02184_));
 sky130_fd_sc_hd__o2111ai_4 _08237_ (.A1(_02172_),
    .A2(_02180_),
    .B1(net29),
    .C1(net63),
    .D1(_02182_),
    .Y(_02185_));
 sky130_fd_sc_hd__o211ai_4 _08238_ (.A1(_00099_),
    .A2(_00396_),
    .B1(_02183_),
    .C1(_02184_),
    .Y(_02186_));
 sky130_fd_sc_hd__o21ai_2 _08239_ (.A1(_02125_),
    .A2(_02126_),
    .B1(_02128_),
    .Y(_02187_));
 sky130_fd_sc_hd__a21oi_4 _08240_ (.A1(_02185_),
    .A2(_02186_),
    .B1(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__and3_1 _08241_ (.A(_02185_),
    .B(_02187_),
    .C(_02186_),
    .X(_02190_));
 sky130_fd_sc_hd__nand3_2 _08242_ (.A(_02185_),
    .B(_02187_),
    .C(_02186_),
    .Y(_02191_));
 sky130_fd_sc_hd__a211o_1 _08243_ (.A1(_02174_),
    .A2(_02177_),
    .B1(_02188_),
    .C1(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__o21ai_2 _08244_ (.A1(_02188_),
    .A2(_02190_),
    .B1(_02179_),
    .Y(_02193_));
 sky130_fd_sc_hd__o21bai_2 _08245_ (.A1(_02188_),
    .A2(_02190_),
    .B1_N(_02179_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand3b_2 _08246_ (.A_N(_02188_),
    .B(_02191_),
    .C(_02179_),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_02194_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(_02192_),
    .B(_02193_),
    .Y(_02197_));
 sky130_fd_sc_hd__o22ai_2 _08249_ (.A1(_02163_),
    .A2(_02168_),
    .B1(_02197_),
    .B2(_02165_),
    .Y(_02198_));
 sky130_fd_sc_hd__a21oi_2 _08250_ (.A1(_02166_),
    .A2(_02196_),
    .B1(_02169_),
    .Y(_02199_));
 sky130_fd_sc_hd__o31a_2 _08251_ (.A1(_00121_),
    .A2(_00385_),
    .A3(_02170_),
    .B1(_02185_),
    .X(_02201_));
 sky130_fd_sc_hd__o21ai_2 _08252_ (.A1(_02170_),
    .A2(_02181_),
    .B1(_02185_),
    .Y(_02202_));
 sky130_fd_sc_hd__o21ai_2 _08253_ (.A1(_02154_),
    .A2(_02155_),
    .B1(_02158_),
    .Y(_02203_));
 sky130_fd_sc_hd__o31a_2 _08254_ (.A1(_00110_),
    .A2(_00352_),
    .A3(_02155_),
    .B1(_02158_),
    .X(_02204_));
 sky130_fd_sc_hd__nand2_2 _08255_ (.A(net32),
    .B(net62),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(net32),
    .B(net61),
    .Y(_02206_));
 sky130_fd_sc_hd__and4_1 _08257_ (.A(net32),
    .B(net31),
    .C(net62),
    .D(net61),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_2 _08258_ (.A1(net31),
    .A2(net62),
    .B1(net61),
    .B2(net32),
    .X(_02208_));
 sky130_fd_sc_hd__o2bb2ai_1 _08259_ (.A1_N(_02180_),
    .A2_N(_02206_),
    .B1(_02205_),
    .B2(_02181_),
    .Y(_02209_));
 sky130_fd_sc_hd__o221ai_4 _08260_ (.A1(_00088_),
    .A2(_00396_),
    .B1(_02181_),
    .B2(_02205_),
    .C1(_02208_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand3_2 _08261_ (.A(_02209_),
    .B(net63),
    .C(net30),
    .Y(_02212_));
 sky130_fd_sc_hd__o21ai_2 _08262_ (.A1(_00088_),
    .A2(_00396_),
    .B1(_02209_),
    .Y(_02213_));
 sky130_fd_sc_hd__o2111ai_4 _08263_ (.A1(_02181_),
    .A2(_02205_),
    .B1(net30),
    .C1(net63),
    .D1(_02208_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand3_4 _08264_ (.A(_02204_),
    .B(_02210_),
    .C(_02212_),
    .Y(_02215_));
 sky130_fd_sc_hd__and3_2 _08265_ (.A(_02213_),
    .B(_02214_),
    .C(_02203_),
    .X(_02216_));
 sky130_fd_sc_hd__nand3_4 _08266_ (.A(_02213_),
    .B(_02214_),
    .C(_02203_),
    .Y(_02217_));
 sky130_fd_sc_hd__a31oi_4 _08267_ (.A1(_02204_),
    .A2(_02210_),
    .A3(_02212_),
    .B1(_02201_),
    .Y(_02218_));
 sky130_fd_sc_hd__and3_2 _08268_ (.A(_02202_),
    .B(_02215_),
    .C(_02217_),
    .X(_02219_));
 sky130_fd_sc_hd__a21oi_4 _08269_ (.A1(_02215_),
    .A2(_02217_),
    .B1(_02202_),
    .Y(_02220_));
 sky130_fd_sc_hd__a21oi_4 _08270_ (.A1(_02215_),
    .A2(_02217_),
    .B1(_02201_),
    .Y(_02221_));
 sky130_fd_sc_hd__and3_2 _08271_ (.A(_02215_),
    .B(_02217_),
    .C(_02201_),
    .X(_02223_));
 sky130_fd_sc_hd__a21o_1 _08272_ (.A1(_02217_),
    .A2(_02218_),
    .B1(_02220_),
    .X(_02224_));
 sky130_fd_sc_hd__a2bb2oi_4 _08273_ (.A1_N(_02151_),
    .A2_N(_02149_),
    .B1(_02161_),
    .B2(_02153_),
    .Y(_02225_));
 sky130_fd_sc_hd__a2bb2o_2 _08274_ (.A1_N(_02151_),
    .A2_N(_02149_),
    .B1(_02161_),
    .B2(_02153_),
    .X(_02226_));
 sky130_fd_sc_hd__o22ai_4 _08275_ (.A1(_02109_),
    .A2(_02141_),
    .B1(_02140_),
    .B2(_02143_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand2_1 _08276_ (.A(net5),
    .B(net55),
    .Y(_02228_));
 sky130_fd_sc_hd__and4_1 _08277_ (.A(net7),
    .B(net6),
    .C(net44),
    .D(net33),
    .X(_02229_));
 sky130_fd_sc_hd__a22oi_2 _08278_ (.A1(net6),
    .A2(net44),
    .B1(net33),
    .B2(net7),
    .Y(_02230_));
 sky130_fd_sc_hd__a22o_1 _08279_ (.A1(net6),
    .A2(net44),
    .B1(net33),
    .B2(net7),
    .X(_02231_));
 sky130_fd_sc_hd__nand3_1 _08280_ (.A(_02141_),
    .B(net33),
    .C(net7),
    .Y(_02232_));
 sky130_fd_sc_hd__nand3_1 _08281_ (.A(_01905_),
    .B(net44),
    .C(net6),
    .Y(_02234_));
 sky130_fd_sc_hd__o2111ai_4 _08282_ (.A1(_01906_),
    .A2(_02142_),
    .B1(net5),
    .C1(net55),
    .D1(_02231_),
    .Y(_02235_));
 sky130_fd_sc_hd__o211ai_4 _08283_ (.A1(_00154_),
    .A2(_00341_),
    .B1(_02232_),
    .C1(_02234_),
    .Y(_02236_));
 sky130_fd_sc_hd__o31a_2 _08284_ (.A1(_02230_),
    .A2(_02228_),
    .A3(_02229_),
    .B1(_02227_),
    .X(_02237_));
 sky130_fd_sc_hd__nand3_2 _08285_ (.A(_02227_),
    .B(_02235_),
    .C(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__a21oi_1 _08286_ (.A1(_02235_),
    .A2(_02236_),
    .B1(_02227_),
    .Y(_02239_));
 sky130_fd_sc_hd__a21o_2 _08287_ (.A1(_02235_),
    .A2(_02236_),
    .B1(_02227_),
    .X(_02240_));
 sky130_fd_sc_hd__nand4_4 _08288_ (.A(net3),
    .B(net4),
    .C(net58),
    .D(net59),
    .Y(_02241_));
 sky130_fd_sc_hd__a22oi_1 _08289_ (.A1(net4),
    .A2(net58),
    .B1(net59),
    .B2(net3),
    .Y(_02242_));
 sky130_fd_sc_hd__a22o_1 _08290_ (.A1(net4),
    .A2(net58),
    .B1(net59),
    .B2(net3),
    .X(_02243_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(net2),
    .B(net60),
    .Y(_02245_));
 sky130_fd_sc_hd__and4_1 _08292_ (.A(_02243_),
    .B(net60),
    .C(net2),
    .D(_02241_),
    .X(_02246_));
 sky130_fd_sc_hd__o2bb2a_1 _08293_ (.A1_N(_02241_),
    .A2_N(_02243_),
    .B1(_00143_),
    .B2(_00352_),
    .X(_02247_));
 sky130_fd_sc_hd__a21o_1 _08294_ (.A1(_02241_),
    .A2(_02243_),
    .B1(_02245_),
    .X(_02248_));
 sky130_fd_sc_hd__o211ai_4 _08295_ (.A1(_00143_),
    .A2(_00352_),
    .B1(_02241_),
    .C1(_02243_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_2 _08296_ (.A(_02248_),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a221oi_4 _08297_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02237_),
    .B2(_02236_),
    .C1(_02239_),
    .Y(_02251_));
 sky130_fd_sc_hd__nand3_1 _08298_ (.A(_02238_),
    .B(_02240_),
    .C(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__a21oi_2 _08299_ (.A1(_02238_),
    .A2(_02240_),
    .B1(_02250_),
    .Y(_02253_));
 sky130_fd_sc_hd__o2bb2ai_2 _08300_ (.A1_N(_02238_),
    .A2_N(_02240_),
    .B1(_02246_),
    .B2(_02247_),
    .Y(_02254_));
 sky130_fd_sc_hd__nand2_1 _08301_ (.A(_02252_),
    .B(_02254_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_2 _08302_ (.A(_02226_),
    .B(_02254_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor3_4 _08303_ (.A(_02225_),
    .B(_02251_),
    .C(_02253_),
    .Y(_02258_));
 sky130_fd_sc_hd__a21oi_4 _08304_ (.A1(_02252_),
    .A2(_02254_),
    .B1(_02226_),
    .Y(_02259_));
 sky130_fd_sc_hd__o21ai_2 _08305_ (.A1(_02251_),
    .A2(_02253_),
    .B1(_02225_),
    .Y(_02260_));
 sky130_fd_sc_hd__o221a_2 _08306_ (.A1(_02221_),
    .A2(_02223_),
    .B1(_02251_),
    .B2(_02257_),
    .C1(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__o221ai_1 _08307_ (.A1(_02221_),
    .A2(_02223_),
    .B1(_02251_),
    .B2(_02257_),
    .C1(_02260_),
    .Y(_02262_));
 sky130_fd_sc_hd__o22ai_2 _08308_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_02258_),
    .B2(_02259_),
    .Y(_02263_));
 sky130_fd_sc_hd__o22ai_4 _08309_ (.A1(_02221_),
    .A2(_02223_),
    .B1(_02258_),
    .B2(_02259_),
    .Y(_02264_));
 sky130_fd_sc_hd__o221ai_4 _08310_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_02251_),
    .B2(_02257_),
    .C1(_02260_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_2 _08311_ (.A(_02263_),
    .B(_02198_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_2 _08312_ (.A1(_02264_),
    .A2(_02265_),
    .B1(_02199_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand3_1 _08313_ (.A(_02263_),
    .B(_02198_),
    .C(_02262_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand3_4 _08314_ (.A(_02199_),
    .B(_02264_),
    .C(_02265_),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_1 _08315_ (.A(net26),
    .B(net36),
    .Y(_02271_));
 sky130_fd_sc_hd__and4_1 _08316_ (.A(net26),
    .B(net23),
    .C(net37),
    .D(net36),
    .X(_02272_));
 sky130_fd_sc_hd__nand4_2 _08317_ (.A(net26),
    .B(net23),
    .C(net37),
    .D(net36),
    .Y(_02273_));
 sky130_fd_sc_hd__a22o_1 _08318_ (.A1(net23),
    .A2(net37),
    .B1(net36),
    .B2(net26),
    .X(_02274_));
 sky130_fd_sc_hd__nand2_1 _08319_ (.A(_02273_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__and4_2 _08320_ (.A(_02274_),
    .B(net38),
    .C(net12),
    .D(_02273_),
    .X(_02276_));
 sky130_fd_sc_hd__a22oi_4 _08321_ (.A1(net12),
    .A2(net38),
    .B1(_02273_),
    .B2(_02274_),
    .Y(_02278_));
 sky130_fd_sc_hd__and3_1 _08322_ (.A(_02275_),
    .B(net38),
    .C(net12),
    .X(_02279_));
 sky130_fd_sc_hd__a21oi_2 _08323_ (.A1(net12),
    .A2(net38),
    .B1(_02275_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _08324_ (.A(_02276_),
    .B(_02278_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_2 _08325_ (.A(net27),
    .B(net34),
    .Y(_02282_));
 sky130_fd_sc_hd__nand4_4 _08326_ (.A(net28),
    .B(net27),
    .C(net64),
    .D(net34),
    .Y(_02283_));
 sky130_fd_sc_hd__a22oi_4 _08327_ (.A1(net28),
    .A2(net64),
    .B1(net34),
    .B2(net27),
    .Y(_02284_));
 sky130_fd_sc_hd__a22o_1 _08328_ (.A1(net28),
    .A2(net64),
    .B1(net34),
    .B2(net27),
    .X(_02285_));
 sky130_fd_sc_hd__nand2_1 _08329_ (.A(net26),
    .B(net35),
    .Y(_02286_));
 sky130_fd_sc_hd__nor3b_2 _08330_ (.A(_02286_),
    .B(_02284_),
    .C_N(_02283_),
    .Y(_02287_));
 sky130_fd_sc_hd__o21ai_4 _08331_ (.A1(_02286_),
    .A2(_02284_),
    .B1(_02283_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand4_4 _08332_ (.A(net28),
    .B(net29),
    .C(net64),
    .D(net34),
    .Y(_02290_));
 sky130_fd_sc_hd__a22oi_1 _08333_ (.A1(net29),
    .A2(net64),
    .B1(net34),
    .B2(net28),
    .Y(_02291_));
 sky130_fd_sc_hd__a22o_1 _08334_ (.A1(net29),
    .A2(net64),
    .B1(net34),
    .B2(net28),
    .X(_02292_));
 sky130_fd_sc_hd__nand3_2 _08335_ (.A(_02292_),
    .B(net27),
    .C(_02290_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand4_2 _08336_ (.A(_02292_),
    .B(net35),
    .C(net27),
    .D(_02290_),
    .Y(_02294_));
 sky130_fd_sc_hd__o2bb2ai_4 _08337_ (.A1_N(_02290_),
    .A2_N(_02292_),
    .B1(_00077_),
    .B2(_00407_),
    .Y(_02295_));
 sky130_fd_sc_hd__o211a_2 _08338_ (.A1(_00407_),
    .A2(_02293_),
    .B1(_02295_),
    .C1(_02289_),
    .X(_02296_));
 sky130_fd_sc_hd__o211ai_4 _08339_ (.A1(_00407_),
    .A2(_02293_),
    .B1(_02295_),
    .C1(_02289_),
    .Y(_02297_));
 sky130_fd_sc_hd__a21oi_2 _08340_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02289_),
    .Y(_02298_));
 sky130_fd_sc_hd__a21o_1 _08341_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02289_),
    .X(_02300_));
 sky130_fd_sc_hd__o22ai_1 _08342_ (.A1(_02276_),
    .A2(_02278_),
    .B1(_02296_),
    .B2(_02298_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand3_1 _08343_ (.A(_02300_),
    .B(_02281_),
    .C(_02297_),
    .Y(_02302_));
 sky130_fd_sc_hd__o211ai_4 _08344_ (.A1(_02276_),
    .A2(_02278_),
    .B1(_02297_),
    .C1(_02300_),
    .Y(_02303_));
 sky130_fd_sc_hd__o22ai_4 _08345_ (.A1(_02279_),
    .A2(_02280_),
    .B1(_02296_),
    .B2(_02298_),
    .Y(_02304_));
 sky130_fd_sc_hd__o21ai_1 _08346_ (.A1(_02179_),
    .A2(_02188_),
    .B1(_02191_),
    .Y(_02305_));
 sky130_fd_sc_hd__o2111ai_4 _08347_ (.A1(_02179_),
    .A2(_02188_),
    .B1(_02191_),
    .C1(_02303_),
    .D1(_02304_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand3_1 _08348_ (.A(_02301_),
    .B(_02302_),
    .C(_02305_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_2 _08349_ (.A(net26),
    .B(net64),
    .Y(_02308_));
 sky130_fd_sc_hd__and4_1 _08350_ (.A(net26),
    .B(net27),
    .C(net64),
    .D(net34),
    .X(_02309_));
 sky130_fd_sc_hd__a22oi_2 _08351_ (.A1(net27),
    .A2(net64),
    .B1(net34),
    .B2(net26),
    .Y(_02311_));
 sky130_fd_sc_hd__a22o_1 _08352_ (.A1(net27),
    .A2(net64),
    .B1(net34),
    .B2(net26),
    .X(_02312_));
 sky130_fd_sc_hd__o2111ai_4 _08353_ (.A1(_02282_),
    .A2(_02308_),
    .B1(net23),
    .C1(net35),
    .D1(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__a31o_1 _08354_ (.A1(_02312_),
    .A2(net35),
    .A3(net23),
    .B1(_02309_),
    .X(_02314_));
 sky130_fd_sc_hd__a22oi_4 _08355_ (.A1(net26),
    .A2(net35),
    .B1(_02283_),
    .B2(_02285_),
    .Y(_02315_));
 sky130_fd_sc_hd__a22o_1 _08356_ (.A1(net26),
    .A2(net35),
    .B1(_02283_),
    .B2(_02285_),
    .X(_02316_));
 sky130_fd_sc_hd__nor2_1 _08357_ (.A(_02287_),
    .B(_02315_),
    .Y(_02317_));
 sky130_fd_sc_hd__o221ai_4 _08358_ (.A1(_02282_),
    .A2(_02308_),
    .B1(_02315_),
    .B2(_02287_),
    .C1(_02313_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand3b_2 _08359_ (.A_N(_02287_),
    .B(_02314_),
    .C(_02316_),
    .Y(_02319_));
 sky130_fd_sc_hd__and4_2 _08360_ (.A(net12),
    .B(net23),
    .C(net37),
    .D(net36),
    .X(_02320_));
 sky130_fd_sc_hd__a22oi_2 _08361_ (.A1(net12),
    .A2(net37),
    .B1(net36),
    .B2(net23),
    .Y(_02322_));
 sky130_fd_sc_hd__a22o_1 _08362_ (.A1(net12),
    .A2(net37),
    .B1(net36),
    .B2(net23),
    .X(_02323_));
 sky130_fd_sc_hd__and4b_1 _08363_ (.A_N(_02320_),
    .B(_02323_),
    .C(net1),
    .D(net38),
    .X(_02324_));
 sky130_fd_sc_hd__o2bb2a_1 _08364_ (.A1_N(net1),
    .A2_N(net38),
    .B1(_02320_),
    .B2(_02322_),
    .X(_02325_));
 sky130_fd_sc_hd__a211oi_2 _08365_ (.A1(net1),
    .A2(net38),
    .B1(_02320_),
    .C1(_02322_),
    .Y(_02326_));
 sky130_fd_sc_hd__o211a_1 _08366_ (.A1(_02320_),
    .A2(_02322_),
    .B1(net1),
    .C1(net38),
    .X(_02327_));
 sky130_fd_sc_hd__o21ai_1 _08367_ (.A1(_02324_),
    .A2(_02325_),
    .B1(_02319_),
    .Y(_02328_));
 sky130_fd_sc_hd__o21a_1 _08368_ (.A1(_02314_),
    .A2(_02317_),
    .B1(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a21oi_2 _08369_ (.A1(_02306_),
    .A2(_02307_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__o2111a_2 _08370_ (.A1(_02314_),
    .A2(_02317_),
    .B1(_02328_),
    .C1(_02307_),
    .D1(_02306_),
    .X(_02331_));
 sky130_fd_sc_hd__nor2_2 _08371_ (.A(_02330_),
    .B(_02331_),
    .Y(_02333_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_02270_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__a21oi_2 _08373_ (.A1(_02270_),
    .A2(_02333_),
    .B1(_02268_),
    .Y(_02335_));
 sky130_fd_sc_hd__o2bb2ai_2 _08374_ (.A1_N(_02333_),
    .A2_N(_02270_),
    .B1(_02267_),
    .B2(_02261_),
    .Y(_02336_));
 sky130_fd_sc_hd__and4_1 _08375_ (.A(net26),
    .B(net27),
    .C(net37),
    .D(net36),
    .X(_02337_));
 sky130_fd_sc_hd__nand4_1 _08376_ (.A(net26),
    .B(net27),
    .C(net37),
    .D(net36),
    .Y(_02338_));
 sky130_fd_sc_hd__a22o_1 _08377_ (.A1(net26),
    .A2(net37),
    .B1(net36),
    .B2(net27),
    .X(_02339_));
 sky130_fd_sc_hd__o21ai_1 _08378_ (.A1(_02026_),
    .A2(_02271_),
    .B1(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__o2111ai_2 _08379_ (.A1(_02026_),
    .A2(_02271_),
    .B1(net23),
    .C1(net38),
    .D1(_02339_),
    .Y(_02341_));
 sky130_fd_sc_hd__a22o_1 _08380_ (.A1(net23),
    .A2(net38),
    .B1(_02338_),
    .B2(_02339_),
    .X(_02342_));
 sky130_fd_sc_hd__a21oi_1 _08381_ (.A1(net23),
    .A2(net38),
    .B1(_02340_),
    .Y(_02344_));
 sky130_fd_sc_hd__and3_1 _08382_ (.A(_02340_),
    .B(net38),
    .C(net23),
    .X(_02345_));
 sky130_fd_sc_hd__nand2_1 _08383_ (.A(_02341_),
    .B(_02342_),
    .Y(_02346_));
 sky130_fd_sc_hd__o31ai_2 _08384_ (.A1(_00077_),
    .A2(_00407_),
    .A3(_02291_),
    .B1(_02290_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _08385_ (.A(net28),
    .B(net35),
    .Y(_02348_));
 sky130_fd_sc_hd__nand4_2 _08386_ (.A(net30),
    .B(net29),
    .C(net64),
    .D(net34),
    .Y(_02349_));
 sky130_fd_sc_hd__a22oi_1 _08387_ (.A1(net30),
    .A2(net64),
    .B1(net34),
    .B2(net29),
    .Y(_02350_));
 sky130_fd_sc_hd__a22o_1 _08388_ (.A1(net30),
    .A2(net64),
    .B1(net34),
    .B2(net29),
    .X(_02351_));
 sky130_fd_sc_hd__o2bb2ai_1 _08389_ (.A1_N(_02349_),
    .A2_N(_02351_),
    .B1(_00066_),
    .B2(_00407_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand4_2 _08390_ (.A(_02351_),
    .B(net35),
    .C(net28),
    .D(_02349_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21oi_1 _08391_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02347_),
    .Y(_02355_));
 sky130_fd_sc_hd__a21o_1 _08392_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02347_),
    .X(_02356_));
 sky130_fd_sc_hd__and3_1 _08393_ (.A(_02347_),
    .B(_02352_),
    .C(_02353_),
    .X(_02357_));
 sky130_fd_sc_hd__nand3_1 _08394_ (.A(_02347_),
    .B(_02352_),
    .C(_02353_),
    .Y(_02358_));
 sky130_fd_sc_hd__o211ai_2 _08395_ (.A1(_02344_),
    .A2(_02345_),
    .B1(_02356_),
    .C1(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__o21ai_2 _08396_ (.A1(_02355_),
    .A2(_02357_),
    .B1(_02346_),
    .Y(_02360_));
 sky130_fd_sc_hd__nand3_1 _08397_ (.A(_02346_),
    .B(_02356_),
    .C(_02358_),
    .Y(_02361_));
 sky130_fd_sc_hd__o22ai_1 _08398_ (.A1(_02344_),
    .A2(_02345_),
    .B1(_02355_),
    .B2(_02357_),
    .Y(_02362_));
 sky130_fd_sc_hd__a21oi_1 _08399_ (.A1(_02202_),
    .A2(_02215_),
    .B1(_02216_),
    .Y(_02363_));
 sky130_fd_sc_hd__o211ai_4 _08400_ (.A1(_02216_),
    .A2(_02218_),
    .B1(_02359_),
    .C1(_02360_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand3_2 _08401_ (.A(_02361_),
    .B(_02362_),
    .C(_02363_),
    .Y(_02366_));
 sky130_fd_sc_hd__o21a_1 _08402_ (.A1(_02279_),
    .A2(_02280_),
    .B1(_02300_),
    .X(_02367_));
 sky130_fd_sc_hd__a31o_1 _08403_ (.A1(_02289_),
    .A2(_02294_),
    .A3(_02295_),
    .B1(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__o211a_2 _08404_ (.A1(_02296_),
    .A2(_02367_),
    .B1(_02366_),
    .C1(_02364_),
    .X(_02369_));
 sky130_fd_sc_hd__o211ai_2 _08405_ (.A1(_02296_),
    .A2(_02367_),
    .B1(_02366_),
    .C1(_02364_),
    .Y(_02370_));
 sky130_fd_sc_hd__a21oi_4 _08406_ (.A1(_02364_),
    .A2(_02366_),
    .B1(_02368_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _08407_ (.A(_02369_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o32a_1 _08408_ (.A1(_02225_),
    .A2(_02251_),
    .A3(_02253_),
    .B1(_02220_),
    .B2(_02219_),
    .X(_02373_));
 sky130_fd_sc_hd__a2bb2oi_2 _08409_ (.A1_N(_02221_),
    .A2_N(_02223_),
    .B1(_02225_),
    .B2(_02256_),
    .Y(_02374_));
 sky130_fd_sc_hd__o22ai_2 _08410_ (.A1(_02251_),
    .A2(_02257_),
    .B1(_02224_),
    .B2(_02259_),
    .Y(_02375_));
 sky130_fd_sc_hd__o21ai_2 _08411_ (.A1(_02245_),
    .A2(_02242_),
    .B1(_02241_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand4_2 _08412_ (.A(net32),
    .B(net2),
    .C(net62),
    .D(net61),
    .Y(_02378_));
 sky130_fd_sc_hd__a22o_1 _08413_ (.A1(net32),
    .A2(net62),
    .B1(net61),
    .B2(net2),
    .X(_02379_));
 sky130_fd_sc_hd__nand3_1 _08414_ (.A(_02205_),
    .B(net61),
    .C(net2),
    .Y(_02380_));
 sky130_fd_sc_hd__nand3_1 _08415_ (.A(_01946_),
    .B(net62),
    .C(net32),
    .Y(_02381_));
 sky130_fd_sc_hd__nand4_4 _08416_ (.A(_02379_),
    .B(net63),
    .C(net31),
    .D(_02378_),
    .Y(_02382_));
 sky130_fd_sc_hd__o211ai_2 _08417_ (.A1(_00121_),
    .A2(_00396_),
    .B1(_02380_),
    .C1(_02381_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand3_2 _08418_ (.A(_02377_),
    .B(_02382_),
    .C(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__a21oi_2 _08419_ (.A1(_02382_),
    .A2(_02383_),
    .B1(_02377_),
    .Y(_02385_));
 sky130_fd_sc_hd__a21o_1 _08420_ (.A1(_02382_),
    .A2(_02383_),
    .B1(_02377_),
    .X(_02386_));
 sky130_fd_sc_hd__a31oi_4 _08421_ (.A1(_02208_),
    .A2(net63),
    .A3(net30),
    .B1(_02207_),
    .Y(_02388_));
 sky130_fd_sc_hd__nor3b_2 _08422_ (.A(_02388_),
    .B(_02385_),
    .C_N(_02384_),
    .Y(_02389_));
 sky130_fd_sc_hd__a21boi_2 _08423_ (.A1(_02384_),
    .A2(_02386_),
    .B1_N(_02388_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_1 _08424_ (.A(_02389_),
    .B(_02390_),
    .Y(_02391_));
 sky130_fd_sc_hd__a22oi_4 _08425_ (.A1(_02236_),
    .A2(_02237_),
    .B1(_02240_),
    .B2(_02250_),
    .Y(_02392_));
 sky130_fd_sc_hd__a22o_1 _08426_ (.A1(_02236_),
    .A2(_02237_),
    .B1(_02240_),
    .B2(_02250_),
    .X(_02393_));
 sky130_fd_sc_hd__o22ai_4 _08427_ (.A1(_01906_),
    .A2(_02142_),
    .B1(_02228_),
    .B2(_02230_),
    .Y(_02394_));
 sky130_fd_sc_hd__o211ai_4 _08428_ (.A1(_00187_),
    .A2(_00341_),
    .B1(_01911_),
    .C1(_01912_),
    .Y(_02395_));
 sky130_fd_sc_hd__o31a_1 _08429_ (.A1(_01908_),
    .A2(_01909_),
    .A3(_01907_),
    .B1(_02394_),
    .X(_02396_));
 sky130_fd_sc_hd__and3_1 _08430_ (.A(_01913_),
    .B(_02394_),
    .C(_02395_),
    .X(_02397_));
 sky130_fd_sc_hd__nand3_2 _08431_ (.A(_01913_),
    .B(_02394_),
    .C(_02395_),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_4 _08432_ (.A1(_01913_),
    .A2(_02395_),
    .B1(_02394_),
    .Y(_02400_));
 sky130_fd_sc_hd__a21o_1 _08433_ (.A1(_01913_),
    .A2(_02395_),
    .B1(_02394_),
    .X(_02401_));
 sky130_fd_sc_hd__a22oi_4 _08434_ (.A1(net5),
    .A2(net58),
    .B1(net59),
    .B2(net4),
    .Y(_02402_));
 sky130_fd_sc_hd__a22o_1 _08435_ (.A1(net5),
    .A2(net58),
    .B1(net59),
    .B2(net4),
    .X(_02403_));
 sky130_fd_sc_hd__and4_1 _08436_ (.A(net5),
    .B(net4),
    .C(net58),
    .D(net59),
    .X(_02404_));
 sky130_fd_sc_hd__nand4_4 _08437_ (.A(net5),
    .B(net4),
    .C(net58),
    .D(net59),
    .Y(_02405_));
 sky130_fd_sc_hd__nand4_1 _08438_ (.A(_02403_),
    .B(_02405_),
    .C(net3),
    .D(net60),
    .Y(_02406_));
 sky130_fd_sc_hd__a22o_1 _08439_ (.A1(net3),
    .A2(net60),
    .B1(_02403_),
    .B2(_02405_),
    .X(_02407_));
 sky130_fd_sc_hd__o211ai_2 _08440_ (.A1(_02402_),
    .A2(_02404_),
    .B1(net3),
    .C1(net60),
    .Y(_02408_));
 sky130_fd_sc_hd__a211o_1 _08441_ (.A1(net3),
    .A2(net60),
    .B1(_02402_),
    .C1(_02404_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_1 _08442_ (.A(_02406_),
    .B(_02407_),
    .Y(_02411_));
 sky130_fd_sc_hd__a221oi_4 _08443_ (.A1(_02408_),
    .A2(_02410_),
    .B1(_02396_),
    .B2(_02395_),
    .C1(_02400_),
    .Y(_02412_));
 sky130_fd_sc_hd__a221o_1 _08444_ (.A1(_02408_),
    .A2(_02410_),
    .B1(_02396_),
    .B2(_02395_),
    .C1(_02400_),
    .X(_02413_));
 sky130_fd_sc_hd__a21boi_4 _08445_ (.A1(_02399_),
    .A2(_02401_),
    .B1_N(_02411_),
    .Y(_02414_));
 sky130_fd_sc_hd__o21ai_1 _08446_ (.A1(_02397_),
    .A2(_02400_),
    .B1(_02411_),
    .Y(_02415_));
 sky130_fd_sc_hd__nor3_4 _08447_ (.A(_02392_),
    .B(_02412_),
    .C(_02414_),
    .Y(_02416_));
 sky130_fd_sc_hd__nand3_4 _08448_ (.A(_02393_),
    .B(_02413_),
    .C(_02415_),
    .Y(_02417_));
 sky130_fd_sc_hd__o21a_1 _08449_ (.A1(_02412_),
    .A2(_02414_),
    .B1(_02392_),
    .X(_02418_));
 sky130_fd_sc_hd__o21ai_4 _08450_ (.A1(_02412_),
    .A2(_02414_),
    .B1(_02392_),
    .Y(_02419_));
 sky130_fd_sc_hd__o211a_1 _08451_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_02417_),
    .C1(_02419_),
    .X(_02421_));
 sky130_fd_sc_hd__o211ai_2 _08452_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_02417_),
    .C1(_02419_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21boi_1 _08453_ (.A1(_02417_),
    .A2(_02419_),
    .B1_N(_02391_),
    .Y(_02423_));
 sky130_fd_sc_hd__o21ai_1 _08454_ (.A1(_02416_),
    .A2(_02418_),
    .B1(_02391_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_2 _08455_ (.A(_02419_),
    .B(_02391_),
    .Y(_02425_));
 sky130_fd_sc_hd__o22ai_2 _08456_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_02416_),
    .B2(_02418_),
    .Y(_02426_));
 sky130_fd_sc_hd__o221a_2 _08457_ (.A1(_02258_),
    .A2(_02374_),
    .B1(_02416_),
    .B2(_02425_),
    .C1(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__o221ai_4 _08458_ (.A1(_02258_),
    .A2(_02374_),
    .B1(_02416_),
    .B2(_02425_),
    .C1(_02426_),
    .Y(_02428_));
 sky130_fd_sc_hd__o211a_1 _08459_ (.A1(_02259_),
    .A2(_02373_),
    .B1(_02422_),
    .C1(_02424_),
    .X(_02429_));
 sky130_fd_sc_hd__o211ai_2 _08460_ (.A1(_02259_),
    .A2(_02373_),
    .B1(_02422_),
    .C1(_02424_),
    .Y(_02430_));
 sky130_fd_sc_hd__o211ai_4 _08461_ (.A1(_02369_),
    .A2(_02371_),
    .B1(_02428_),
    .C1(_02430_),
    .Y(_02432_));
 sky130_fd_sc_hd__o21ai_2 _08462_ (.A1(_02427_),
    .A2(_02429_),
    .B1(_02372_),
    .Y(_02433_));
 sky130_fd_sc_hd__o31ai_2 _08463_ (.A1(_02375_),
    .A2(_02421_),
    .A3(_02423_),
    .B1(_02372_),
    .Y(_02434_));
 sky130_fd_sc_hd__o22ai_2 _08464_ (.A1(_02369_),
    .A2(_02371_),
    .B1(_02427_),
    .B2(_02429_),
    .Y(_02435_));
 sky130_fd_sc_hd__o211a_1 _08465_ (.A1(_02434_),
    .A2(_02427_),
    .B1(_02336_),
    .C1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__o211ai_4 _08466_ (.A1(_02434_),
    .A2(_02427_),
    .B1(_02336_),
    .C1(_02435_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21boi_2 _08467_ (.A1(_02306_),
    .A2(_02329_),
    .B1_N(_02307_),
    .Y(_02438_));
 sky130_fd_sc_hd__a31o_1 _08468_ (.A1(_02323_),
    .A2(net38),
    .A3(net1),
    .B1(_02320_),
    .X(_02439_));
 sky130_fd_sc_hd__and3_1 _08469_ (.A(_02439_),
    .B(net39),
    .C(net1),
    .X(_02440_));
 sky130_fd_sc_hd__or3b_4 _08470_ (.A(_00033_),
    .B(_00440_),
    .C_N(_02439_),
    .X(_02441_));
 sky130_fd_sc_hd__nand4_4 _08471_ (.A(net12),
    .B(net1),
    .C(net39),
    .D(net40),
    .Y(_02443_));
 sky130_fd_sc_hd__a22o_1 _08472_ (.A1(net12),
    .A2(net39),
    .B1(net40),
    .B2(net1),
    .X(_02444_));
 sky130_fd_sc_hd__o211ai_4 _08473_ (.A1(_02272_),
    .A2(_02276_),
    .B1(_02443_),
    .C1(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__a211o_1 _08474_ (.A1(_02443_),
    .A2(_02444_),
    .B1(_02272_),
    .C1(_02276_),
    .X(_02446_));
 sky130_fd_sc_hd__nand2_1 _08475_ (.A(_02445_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__and3_2 _08476_ (.A(_02446_),
    .B(_02440_),
    .C(_02445_),
    .X(_02448_));
 sky130_fd_sc_hd__a21oi_1 _08477_ (.A1(_02445_),
    .A2(_02446_),
    .B1(_02440_),
    .Y(_02449_));
 sky130_fd_sc_hd__or2_1 _08478_ (.A(_02448_),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__nor2_1 _08479_ (.A(_02438_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__or3_1 _08480_ (.A(_02438_),
    .B(_02448_),
    .C(_02449_),
    .X(_02452_));
 sky130_fd_sc_hd__o21ai_2 _08481_ (.A1(_02448_),
    .A2(_02449_),
    .B1(_02438_),
    .Y(_02454_));
 sky130_fd_sc_hd__and2b_1 _08482_ (.A_N(_02451_),
    .B(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__nand2b_1 _08483_ (.A_N(_02451_),
    .B(_02454_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand3_1 _08484_ (.A(_02433_),
    .B(_02335_),
    .C(_02432_),
    .Y(_02457_));
 sky130_fd_sc_hd__a31oi_4 _08485_ (.A1(_02433_),
    .A2(_02335_),
    .A3(_02432_),
    .B1(_02456_),
    .Y(_02458_));
 sky130_fd_sc_hd__a31o_1 _08486_ (.A1(_02433_),
    .A2(_02335_),
    .A3(_02432_),
    .B1(_02456_),
    .X(_02459_));
 sky130_fd_sc_hd__and3_1 _08487_ (.A(_02437_),
    .B(_02457_),
    .C(_02455_),
    .X(_02460_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_02458_),
    .B(_02437_),
    .Y(_02461_));
 sky130_fd_sc_hd__a21o_1 _08489_ (.A1(_02457_),
    .A2(_02455_),
    .B1(_02436_),
    .X(_02462_));
 sky130_fd_sc_hd__o21a_1 _08490_ (.A1(_02388_),
    .A2(_02385_),
    .B1(_02384_),
    .X(_02463_));
 sky130_fd_sc_hd__o21ai_2 _08491_ (.A1(_02388_),
    .A2(_02385_),
    .B1(_02384_),
    .Y(_02465_));
 sky130_fd_sc_hd__a22oi_4 _08492_ (.A1(net26),
    .A2(net38),
    .B1(_02028_),
    .B2(_02029_),
    .Y(_02466_));
 sky130_fd_sc_hd__and4_2 _08493_ (.A(_02028_),
    .B(_02029_),
    .C(net26),
    .D(net38),
    .X(_02467_));
 sky130_fd_sc_hd__nor2_2 _08494_ (.A(_02466_),
    .B(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__o211ai_2 _08495_ (.A1(_00099_),
    .A2(_00407_),
    .B1(_01992_),
    .C1(_01993_),
    .Y(_02469_));
 sky130_fd_sc_hd__o21ai_2 _08496_ (.A1(_02348_),
    .A2(_02350_),
    .B1(_02349_),
    .Y(_02470_));
 sky130_fd_sc_hd__and3_2 _08497_ (.A(_01994_),
    .B(_02470_),
    .C(_02469_),
    .X(_02471_));
 sky130_fd_sc_hd__nand3_2 _08498_ (.A(_01994_),
    .B(_02470_),
    .C(_02469_),
    .Y(_02472_));
 sky130_fd_sc_hd__a21oi_1 _08499_ (.A1(_01994_),
    .A2(_02469_),
    .B1(_02470_),
    .Y(_02473_));
 sky130_fd_sc_hd__a21o_2 _08500_ (.A1(_01994_),
    .A2(_02469_),
    .B1(_02470_),
    .X(_02474_));
 sky130_fd_sc_hd__o21ai_2 _08501_ (.A1(_02471_),
    .A2(_02473_),
    .B1(_02468_),
    .Y(_02476_));
 sky130_fd_sc_hd__o211ai_4 _08502_ (.A1(_02466_),
    .A2(_02467_),
    .B1(_02472_),
    .C1(_02474_),
    .Y(_02477_));
 sky130_fd_sc_hd__o22ai_1 _08503_ (.A1(_02466_),
    .A2(_02467_),
    .B1(_02471_),
    .B2(_02473_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand3_1 _08504_ (.A(_02468_),
    .B(_02472_),
    .C(_02474_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand3_2 _08505_ (.A(_02476_),
    .B(_02477_),
    .C(_02463_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand3_2 _08506_ (.A(_02465_),
    .B(_02478_),
    .C(_02479_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21o_1 _08507_ (.A1(_02346_),
    .A2(_02358_),
    .B1(_02355_),
    .X(_02482_));
 sky130_fd_sc_hd__a31o_1 _08508_ (.A1(_02341_),
    .A2(_02342_),
    .A3(_02356_),
    .B1(_02357_),
    .X(_02483_));
 sky130_fd_sc_hd__a21oi_2 _08509_ (.A1(_02480_),
    .A2(_02481_),
    .B1(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__a21o_1 _08510_ (.A1(_02480_),
    .A2(_02481_),
    .B1(_02483_),
    .X(_02485_));
 sky130_fd_sc_hd__and3_1 _08511_ (.A(_02480_),
    .B(_02481_),
    .C(_02483_),
    .X(_02487_));
 sky130_fd_sc_hd__nand3_1 _08512_ (.A(_02480_),
    .B(_02481_),
    .C(_02483_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _08513_ (.A(_02484_),
    .B(_02487_),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(_02485_),
    .B(_02488_),
    .Y(_02490_));
 sky130_fd_sc_hd__a21oi_1 _08515_ (.A1(_02419_),
    .A2(_02391_),
    .B1(_02416_),
    .Y(_02491_));
 sky130_fd_sc_hd__a21o_1 _08516_ (.A1(_02419_),
    .A2(_02391_),
    .B1(_02416_),
    .X(_02492_));
 sky130_fd_sc_hd__o31a_2 _08517_ (.A1(_00110_),
    .A2(_00374_),
    .A3(_01946_),
    .B1(_02382_),
    .X(_02493_));
 sky130_fd_sc_hd__o31a_1 _08518_ (.A1(_00132_),
    .A2(_00352_),
    .A3(_02402_),
    .B1(_02405_),
    .X(_02494_));
 sky130_fd_sc_hd__o31ai_4 _08519_ (.A1(_00132_),
    .A2(_00352_),
    .A3(_02402_),
    .B1(_02405_),
    .Y(_02495_));
 sky130_fd_sc_hd__o2bb2ai_2 _08520_ (.A1_N(_01949_),
    .A2_N(_01950_),
    .B1(_00110_),
    .B2(_00396_),
    .Y(_02496_));
 sky130_fd_sc_hd__nand2_1 _08521_ (.A(_01952_),
    .B(_02496_),
    .Y(_02498_));
 sky130_fd_sc_hd__a21oi_2 _08522_ (.A1(_01952_),
    .A2(_02496_),
    .B1(_02495_),
    .Y(_02499_));
 sky130_fd_sc_hd__a21o_1 _08523_ (.A1(_01952_),
    .A2(_02496_),
    .B1(_02495_),
    .X(_02500_));
 sky130_fd_sc_hd__and3_2 _08524_ (.A(_01952_),
    .B(_02495_),
    .C(_02496_),
    .X(_02501_));
 sky130_fd_sc_hd__nand3_2 _08525_ (.A(_01952_),
    .B(_02495_),
    .C(_02496_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand3b_4 _08526_ (.A_N(_02493_),
    .B(_02500_),
    .C(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__o21ai_4 _08527_ (.A1(_02499_),
    .A2(_02501_),
    .B1(_02493_),
    .Y(_02504_));
 sky130_fd_sc_hd__a22o_1 _08528_ (.A1(_02378_),
    .A2(_02382_),
    .B1(_02500_),
    .B2(_02502_),
    .X(_02505_));
 sky130_fd_sc_hd__nand4_1 _08529_ (.A(_02378_),
    .B(_02382_),
    .C(_02500_),
    .D(_02502_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2_1 _08530_ (.A(_02505_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _08531_ (.A(_02503_),
    .B(_02504_),
    .Y(_02509_));
 sky130_fd_sc_hd__o2bb2a_1 _08532_ (.A1_N(_02395_),
    .A2_N(_02396_),
    .B1(_02400_),
    .B2(_02411_),
    .X(_02510_));
 sky130_fd_sc_hd__o21ai_2 _08533_ (.A1(_02400_),
    .A2(_02411_),
    .B1(_02399_),
    .Y(_02511_));
 sky130_fd_sc_hd__a21boi_2 _08534_ (.A1(_01920_),
    .A2(_01922_),
    .B1_N(_01934_),
    .Y(_02512_));
 sky130_fd_sc_hd__o2bb2ai_4 _08535_ (.A1_N(_01920_),
    .A2_N(_01922_),
    .B1(_01930_),
    .B2(_01932_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _08536_ (.A(_01937_),
    .B(_02513_),
    .Y(_02514_));
 sky130_fd_sc_hd__a21oi_1 _08537_ (.A1(_01937_),
    .A2(_02513_),
    .B1(_02511_),
    .Y(_02515_));
 sky130_fd_sc_hd__o21ai_4 _08538_ (.A1(_01935_),
    .A2(_02512_),
    .B1(_02510_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand2_2 _08539_ (.A(_02511_),
    .B(_02513_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand3_4 _08540_ (.A(_01937_),
    .B(_02511_),
    .C(_02513_),
    .Y(_02518_));
 sky130_fd_sc_hd__a22oi_4 _08541_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_02516_),
    .B2(_02518_),
    .Y(_02520_));
 sky130_fd_sc_hd__a22o_1 _08542_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_02516_),
    .B2(_02518_),
    .X(_02521_));
 sky130_fd_sc_hd__a22oi_2 _08543_ (.A1(_02505_),
    .A2(_02506_),
    .B1(_02514_),
    .B2(_02510_),
    .Y(_02522_));
 sky130_fd_sc_hd__o211a_1 _08544_ (.A1(_01935_),
    .A2(_02517_),
    .B1(_02516_),
    .C1(_02507_),
    .X(_02523_));
 sky130_fd_sc_hd__o2111ai_4 _08545_ (.A1(_01935_),
    .A2(_02517_),
    .B1(_02516_),
    .C1(_02504_),
    .D1(_02503_),
    .Y(_02524_));
 sky130_fd_sc_hd__a221oi_4 _08546_ (.A1(_02522_),
    .A2(_02518_),
    .B1(_02425_),
    .B2(_02417_),
    .C1(_02520_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand3_2 _08547_ (.A(_02492_),
    .B(_02521_),
    .C(_02524_),
    .Y(_02526_));
 sky130_fd_sc_hd__a21oi_2 _08548_ (.A1(_02521_),
    .A2(_02524_),
    .B1(_02492_),
    .Y(_02527_));
 sky130_fd_sc_hd__o21ai_2 _08549_ (.A1(_02520_),
    .A2(_02523_),
    .B1(_02491_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand4_4 _08550_ (.A(_02485_),
    .B(_02488_),
    .C(_02526_),
    .D(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__o22ai_4 _08551_ (.A1(_02484_),
    .A2(_02487_),
    .B1(_02525_),
    .B2(_02527_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _08552_ (.A(_02529_),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21a_1 _08553_ (.A1(_02369_),
    .A2(_02371_),
    .B1(_02428_),
    .X(_02533_));
 sky130_fd_sc_hd__o32a_1 _08554_ (.A1(_02375_),
    .A2(_02421_),
    .A3(_02423_),
    .B1(_02427_),
    .B2(_02372_),
    .X(_02534_));
 sky130_fd_sc_hd__o31a_1 _08555_ (.A1(_02369_),
    .A2(_02371_),
    .A3(_02429_),
    .B1(_02428_),
    .X(_02535_));
 sky130_fd_sc_hd__nand3_2 _08556_ (.A(_02534_),
    .B(_02531_),
    .C(_02529_),
    .Y(_02536_));
 sky130_fd_sc_hd__a21oi_1 _08557_ (.A1(_02529_),
    .A2(_02531_),
    .B1(_02534_),
    .Y(_02537_));
 sky130_fd_sc_hd__o2bb2ai_2 _08558_ (.A1_N(_02529_),
    .A2_N(_02531_),
    .B1(_02533_),
    .B2(_02429_),
    .Y(_02538_));
 sky130_fd_sc_hd__a31o_1 _08559_ (.A1(_02339_),
    .A2(net38),
    .A3(net23),
    .B1(_02337_),
    .X(_02539_));
 sky130_fd_sc_hd__o22ai_2 _08560_ (.A1(_00033_),
    .A2(_00451_),
    .B1(_02040_),
    .B2(_02041_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21oi_1 _08561_ (.A1(_02044_),
    .A2(_02540_),
    .B1(_02539_),
    .Y(_02542_));
 sky130_fd_sc_hd__a21o_1 _08562_ (.A1(_02044_),
    .A2(_02540_),
    .B1(_02539_),
    .X(_02543_));
 sky130_fd_sc_hd__nand3_1 _08563_ (.A(_02044_),
    .B(_02539_),
    .C(_02540_),
    .Y(_02544_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(_02543_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand3_1 _08565_ (.A(_02443_),
    .B(_02445_),
    .C(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _08566_ (.A1(_02443_),
    .A2(_02445_),
    .B1(_02545_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _08567_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__and3_1 _08568_ (.A(_02364_),
    .B(_02370_),
    .C(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__nand3_1 _08569_ (.A(_02364_),
    .B(_02370_),
    .C(_02548_),
    .Y(_02550_));
 sky130_fd_sc_hd__a21oi_2 _08570_ (.A1(_02364_),
    .A2(_02370_),
    .B1(_02548_),
    .Y(_02551_));
 sky130_fd_sc_hd__o22a_1 _08571_ (.A1(_02441_),
    .A2(_02447_),
    .B1(_02549_),
    .B2(_02551_),
    .X(_02553_));
 sky130_fd_sc_hd__o22ai_2 _08572_ (.A1(_02441_),
    .A2(_02447_),
    .B1(_02549_),
    .B2(_02551_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor4_1 _08573_ (.A(_02441_),
    .B(_02447_),
    .C(_02549_),
    .D(_02551_),
    .Y(_02555_));
 sky130_fd_sc_hd__nand3b_2 _08574_ (.A_N(_02551_),
    .B(_02448_),
    .C(_02550_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _08575_ (.A(_02554_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__nand4_4 _08576_ (.A(_02536_),
    .B(_02538_),
    .C(_02554_),
    .D(_02556_),
    .Y(_02558_));
 sky130_fd_sc_hd__o2bb2ai_2 _08577_ (.A1_N(_02536_),
    .A2_N(_02538_),
    .B1(_02553_),
    .B2(_02555_),
    .Y(_02559_));
 sky130_fd_sc_hd__o211a_1 _08578_ (.A1(_02436_),
    .A2(_02458_),
    .B1(_02558_),
    .C1(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__o211ai_1 _08579_ (.A1(_02436_),
    .A2(_02458_),
    .B1(_02558_),
    .C1(_02559_),
    .Y(_02561_));
 sky130_fd_sc_hd__a21oi_1 _08580_ (.A1(_02558_),
    .A2(_02559_),
    .B1(_02462_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21o_1 _08581_ (.A1(_02558_),
    .A2(_02559_),
    .B1(_02462_),
    .X(_02564_));
 sky130_fd_sc_hd__nand3b_1 _08582_ (.A_N(_02452_),
    .B(_02561_),
    .C(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__o31a_1 _08583_ (.A1(_02438_),
    .A2(_02450_),
    .A3(_02562_),
    .B1(_02561_),
    .X(_02566_));
 sky130_fd_sc_hd__o21ai_1 _08584_ (.A1(_02557_),
    .A2(_02537_),
    .B1(_02536_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(_02445_),
    .B(_02545_),
    .Y(_02568_));
 sky130_fd_sc_hd__a21oi_2 _08586_ (.A1(_02038_),
    .A2(_02047_),
    .B1(_02045_),
    .Y(_02569_));
 sky130_fd_sc_hd__a21o_1 _08587_ (.A1(_02038_),
    .A2(_02047_),
    .B1(_02045_),
    .X(_02570_));
 sky130_fd_sc_hd__o21ai_2 _08588_ (.A1(_02443_),
    .A2(_02542_),
    .B1(_02544_),
    .Y(_02571_));
 sky130_fd_sc_hd__o21a_1 _08589_ (.A1(_02443_),
    .A2(_02542_),
    .B1(_02544_),
    .X(_02572_));
 sky130_fd_sc_hd__o21ai_4 _08590_ (.A1(_02049_),
    .A2(_02569_),
    .B1(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__inv_2 _08591_ (.A(_02573_),
    .Y(_02575_));
 sky130_fd_sc_hd__o211ai_4 _08592_ (.A1(_02037_),
    .A2(_02048_),
    .B1(_02571_),
    .C1(_02570_),
    .Y(_02576_));
 sky130_fd_sc_hd__o211ai_1 _08593_ (.A1(_00033_),
    .A2(_00473_),
    .B1(_02573_),
    .C1(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21o_1 _08594_ (.A1(_02573_),
    .A2(_02576_),
    .B1(_01851_),
    .X(_02578_));
 sky130_fd_sc_hd__o2bb2ai_1 _08595_ (.A1_N(_02573_),
    .A2_N(_02576_),
    .B1(_00033_),
    .B2(_00473_),
    .Y(_02579_));
 sky130_fd_sc_hd__and4_1 _08596_ (.A(_02573_),
    .B(_02576_),
    .C(net1),
    .D(net42),
    .X(_02580_));
 sky130_fd_sc_hd__nand4_1 _08597_ (.A(_02573_),
    .B(_02576_),
    .C(net1),
    .D(net42),
    .Y(_02581_));
 sky130_fd_sc_hd__a32oi_2 _08598_ (.A1(_02463_),
    .A2(_02476_),
    .A3(_02477_),
    .B1(_02481_),
    .B2(_02482_),
    .Y(_02582_));
 sky130_fd_sc_hd__a32o_1 _08599_ (.A1(_02463_),
    .A2(_02476_),
    .A3(_02477_),
    .B1(_02481_),
    .B2(_02482_),
    .X(_02583_));
 sky130_fd_sc_hd__nand3_2 _08600_ (.A(_02577_),
    .B(_02578_),
    .C(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _08601_ (.A(_02579_),
    .B(_02582_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand3_1 _08602_ (.A(_02579_),
    .B(_02581_),
    .C(_02582_),
    .Y(_02587_));
 sky130_fd_sc_hd__a21oi_1 _08603_ (.A1(_02584_),
    .A2(_02587_),
    .B1(_02568_),
    .Y(_02588_));
 sky130_fd_sc_hd__a2bb2o_1 _08604_ (.A1_N(_02445_),
    .A2_N(_02545_),
    .B1(_02584_),
    .B2(_02587_),
    .X(_02589_));
 sky130_fd_sc_hd__and3_1 _08605_ (.A(_02584_),
    .B(_02587_),
    .C(_02568_),
    .X(_02590_));
 sky130_fd_sc_hd__o211ai_1 _08606_ (.A1(_02580_),
    .A2(_02586_),
    .B1(_02584_),
    .C1(_02568_),
    .Y(_02591_));
 sky130_fd_sc_hd__nor2_1 _08607_ (.A(_02588_),
    .B(_02590_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _08608_ (.A1(_02528_),
    .A2(_02489_),
    .B1(_02525_),
    .Y(_02593_));
 sky130_fd_sc_hd__o21ai_1 _08609_ (.A1(_02490_),
    .A2(_02527_),
    .B1(_02526_),
    .Y(_02594_));
 sky130_fd_sc_hd__o2bb2a_1 _08610_ (.A1_N(_01998_),
    .A2_N(_02000_),
    .B1(_02001_),
    .B2(_01828_),
    .X(_02595_));
 sky130_fd_sc_hd__o2bb2ai_2 _08611_ (.A1_N(_01998_),
    .A2_N(_02000_),
    .B1(_02001_),
    .B2(_01828_),
    .Y(_02597_));
 sky130_fd_sc_hd__nand3b_2 _08612_ (.A_N(_02004_),
    .B(_02000_),
    .C(_01998_),
    .Y(_02598_));
 sky130_fd_sc_hd__a21oi_2 _08613_ (.A1(_02498_),
    .A2(_02494_),
    .B1(_02493_),
    .Y(_02599_));
 sky130_fd_sc_hd__o21ai_1 _08614_ (.A1(_02493_),
    .A2(_02499_),
    .B1(_02502_),
    .Y(_02600_));
 sky130_fd_sc_hd__a21oi_1 _08615_ (.A1(_02597_),
    .A2(_02598_),
    .B1(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__a21o_1 _08616_ (.A1(_02597_),
    .A2(_02598_),
    .B1(_02600_),
    .X(_02602_));
 sky130_fd_sc_hd__o21ai_1 _08617_ (.A1(_02501_),
    .A2(_02599_),
    .B1(_02598_),
    .Y(_02603_));
 sky130_fd_sc_hd__o211a_1 _08618_ (.A1(_02501_),
    .A2(_02599_),
    .B1(_02598_),
    .C1(_02597_),
    .X(_02604_));
 sky130_fd_sc_hd__o211ai_2 _08619_ (.A1(_02501_),
    .A2(_02599_),
    .B1(_02598_),
    .C1(_02597_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21ai_2 _08620_ (.A1(_02468_),
    .A2(_02471_),
    .B1(_02474_),
    .Y(_02606_));
 sky130_fd_sc_hd__o2111ai_4 _08621_ (.A1(_02468_),
    .A2(_02471_),
    .B1(_02474_),
    .C1(_02602_),
    .D1(_02605_),
    .Y(_02608_));
 sky130_fd_sc_hd__o21ai_2 _08622_ (.A1(_02601_),
    .A2(_02604_),
    .B1(_02606_),
    .Y(_02609_));
 sky130_fd_sc_hd__nand2_2 _08623_ (.A(_02608_),
    .B(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hd__o2bb2ai_4 _08624_ (.A1_N(_01944_),
    .A2_N(_01945_),
    .B1(_01960_),
    .B2(_01961_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand3_2 _08625_ (.A(_01944_),
    .B(_01945_),
    .C(_01962_),
    .Y(_02612_));
 sky130_fd_sc_hd__o22ai_4 _08626_ (.A1(_01935_),
    .A2(_02517_),
    .B1(_02509_),
    .B2(_02515_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_4 _08627_ (.A1(_02611_),
    .A2(_02612_),
    .B1(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a21o_1 _08628_ (.A1(_02611_),
    .A2(_02612_),
    .B1(_02613_),
    .X(_02615_));
 sky130_fd_sc_hd__o211a_1 _08629_ (.A1(_01943_),
    .A2(_01963_),
    .B1(_02611_),
    .C1(_02613_),
    .X(_02616_));
 sky130_fd_sc_hd__o211ai_4 _08630_ (.A1(_01943_),
    .A2(_01963_),
    .B1(_02611_),
    .C1(_02613_),
    .Y(_02617_));
 sky130_fd_sc_hd__o21bai_2 _08631_ (.A1(_02614_),
    .A2(_02616_),
    .B1_N(_02610_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand3_1 _08632_ (.A(_02610_),
    .B(_02615_),
    .C(_02617_),
    .Y(_02620_));
 sky130_fd_sc_hd__nand4_1 _08633_ (.A(_02608_),
    .B(_02609_),
    .C(_02615_),
    .D(_02617_),
    .Y(_02621_));
 sky130_fd_sc_hd__o21ai_1 _08634_ (.A1(_02614_),
    .A2(_02616_),
    .B1(_02610_),
    .Y(_02622_));
 sky130_fd_sc_hd__a21oi_1 _08635_ (.A1(_02619_),
    .A2(_02620_),
    .B1(_02593_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand3_1 _08636_ (.A(_02594_),
    .B(_02621_),
    .C(_02622_),
    .Y(_02624_));
 sky130_fd_sc_hd__o2111a_1 _08637_ (.A1(_02527_),
    .A2(_02490_),
    .B1(_02526_),
    .C1(_02619_),
    .D1(_02620_),
    .X(_02625_));
 sky130_fd_sc_hd__nand3_2 _08638_ (.A(_02593_),
    .B(_02619_),
    .C(_02620_),
    .Y(_02626_));
 sky130_fd_sc_hd__o211ai_1 _08639_ (.A1(_02588_),
    .A2(_02590_),
    .B1(_02624_),
    .C1(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__o21ai_1 _08640_ (.A1(_02623_),
    .A2(_02625_),
    .B1(_02592_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand4_1 _08641_ (.A(_02589_),
    .B(_02591_),
    .C(_02624_),
    .D(_02626_),
    .Y(_02630_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(_02589_),
    .A2(_02591_),
    .B1(_02624_),
    .B2(_02626_),
    .X(_02631_));
 sky130_fd_sc_hd__o2111ai_2 _08643_ (.A1(_02532_),
    .A2(_02535_),
    .B1(_02558_),
    .C1(_02627_),
    .D1(_02628_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand3_1 _08644_ (.A(_02567_),
    .B(_02630_),
    .C(_02631_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21oi_1 _08645_ (.A1(_02448_),
    .A2(_02550_),
    .B1(_02551_),
    .Y(_02634_));
 sky130_fd_sc_hd__a21oi_1 _08646_ (.A1(_02632_),
    .A2(_02633_),
    .B1(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__and3_1 _08647_ (.A(_02632_),
    .B(_02633_),
    .C(_02634_),
    .X(_02636_));
 sky130_fd_sc_hd__nor2_1 _08648_ (.A(_02635_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__o22ai_1 _08649_ (.A1(_02438_),
    .A2(_02450_),
    .B1(_02560_),
    .B2(_02562_),
    .Y(_02638_));
 sky130_fd_sc_hd__nand2_1 _08650_ (.A(net2),
    .B(net44),
    .Y(_02639_));
 sky130_fd_sc_hd__a22oi_2 _08651_ (.A1(net2),
    .A2(net44),
    .B1(net33),
    .B2(net3),
    .Y(_02641_));
 sky130_fd_sc_hd__a22o_2 _08652_ (.A1(net2),
    .A2(net44),
    .B1(net33),
    .B2(net3),
    .X(_02642_));
 sky130_fd_sc_hd__and4_2 _08653_ (.A(net3),
    .B(net2),
    .C(net44),
    .D(net33),
    .X(_02643_));
 sky130_fd_sc_hd__nand4_1 _08654_ (.A(net3),
    .B(net2),
    .C(net44),
    .D(net33),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(net32),
    .B(net55),
    .Y(_02645_));
 sky130_fd_sc_hd__o21ai_2 _08656_ (.A1(_02096_),
    .A2(_02639_),
    .B1(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__a21oi_1 _08657_ (.A1(_02096_),
    .A2(_02639_),
    .B1(_02645_),
    .Y(_02647_));
 sky130_fd_sc_hd__and3_1 _08658_ (.A(_02100_),
    .B(_02104_),
    .C(_02105_),
    .X(_02648_));
 sky130_fd_sc_hd__o211ai_4 _08659_ (.A1(_00143_),
    .A2(_00341_),
    .B1(_02104_),
    .C1(_02105_),
    .Y(_02649_));
 sky130_fd_sc_hd__o21ai_2 _08660_ (.A1(_02643_),
    .A2(_02647_),
    .B1(_02106_),
    .Y(_02650_));
 sky130_fd_sc_hd__o211a_2 _08661_ (.A1(_02643_),
    .A2(_02647_),
    .B1(_02649_),
    .C1(_02106_),
    .X(_02652_));
 sky130_fd_sc_hd__and4_1 _08662_ (.A(net32),
    .B(net31),
    .C(net58),
    .D(net59),
    .X(_02653_));
 sky130_fd_sc_hd__nand4_2 _08663_ (.A(net32),
    .B(net31),
    .C(net58),
    .D(net59),
    .Y(_02654_));
 sky130_fd_sc_hd__a22o_1 _08664_ (.A1(net32),
    .A2(net58),
    .B1(net59),
    .B2(net31),
    .X(_02655_));
 sky130_fd_sc_hd__o2bb2a_1 _08665_ (.A1_N(_02654_),
    .A2_N(_02655_),
    .B1(_00088_),
    .B2(_00352_),
    .X(_02656_));
 sky130_fd_sc_hd__a22o_1 _08666_ (.A1(net30),
    .A2(net60),
    .B1(_02654_),
    .B2(_02655_),
    .X(_02657_));
 sky130_fd_sc_hd__and4_2 _08667_ (.A(_02655_),
    .B(net60),
    .C(net30),
    .D(_02654_),
    .X(_02658_));
 sky130_fd_sc_hd__nand4_2 _08668_ (.A(_02655_),
    .B(net60),
    .C(net30),
    .D(_02654_),
    .Y(_02659_));
 sky130_fd_sc_hd__a22oi_4 _08669_ (.A1(_02642_),
    .A2(_02646_),
    .B1(_02649_),
    .B2(_02106_),
    .Y(_02660_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(_02642_),
    .A2(_02646_),
    .B1(_02649_),
    .B2(_02106_),
    .X(_02661_));
 sky130_fd_sc_hd__o2111a_2 _08671_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_02657_),
    .C1(_02659_),
    .D1(_02661_),
    .X(_02663_));
 sky130_fd_sc_hd__o2111ai_4 _08672_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_02657_),
    .C1(_02659_),
    .D1(_02661_),
    .Y(_02664_));
 sky130_fd_sc_hd__o32a_2 _08673_ (.A1(_02656_),
    .A2(_02658_),
    .A3(_02660_),
    .B1(_02650_),
    .B2(_02648_),
    .X(_02665_));
 sky130_fd_sc_hd__a31o_1 _08674_ (.A1(_02657_),
    .A2(_02659_),
    .A3(_02661_),
    .B1(_02652_),
    .X(_02666_));
 sky130_fd_sc_hd__a21oi_1 _08675_ (.A1(_02121_),
    .A2(_02124_),
    .B1(_02135_),
    .Y(_02667_));
 sky130_fd_sc_hd__o2bb2ai_2 _08676_ (.A1_N(_02121_),
    .A2_N(_02124_),
    .B1(_02131_),
    .B2(_02132_),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _08677_ (.A(_02137_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__o211ai_4 _08678_ (.A1(_02652_),
    .A2(_02663_),
    .B1(_02668_),
    .C1(_02137_),
    .Y(_02670_));
 sky130_fd_sc_hd__a21oi_1 _08679_ (.A1(_02137_),
    .A2(_02668_),
    .B1(_02666_),
    .Y(_02671_));
 sky130_fd_sc_hd__o21ai_4 _08680_ (.A1(_02136_),
    .A2(_02667_),
    .B1(_02665_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_1 _08681_ (.A(net28),
    .B(net61),
    .Y(_02674_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(net28),
    .B(net62),
    .Y(_02675_));
 sky130_fd_sc_hd__and2_1 _08683_ (.A(net27),
    .B(net63),
    .X(_02676_));
 sky130_fd_sc_hd__a22o_1 _08684_ (.A1(net28),
    .A2(net62),
    .B1(net61),
    .B2(net29),
    .X(_02677_));
 sky130_fd_sc_hd__nand3_1 _08685_ (.A(_02675_),
    .B(net61),
    .C(net29),
    .Y(_02678_));
 sky130_fd_sc_hd__nand3_1 _08686_ (.A(_02171_),
    .B(net62),
    .C(net28),
    .Y(_02679_));
 sky130_fd_sc_hd__o211ai_2 _08687_ (.A1(_02173_),
    .A2(_02674_),
    .B1(_02676_),
    .C1(_02677_),
    .Y(_02680_));
 sky130_fd_sc_hd__a2bb2o_2 _08688_ (.A1_N(_02173_),
    .A2_N(_02674_),
    .B1(_02676_),
    .B2(_02677_),
    .X(_02681_));
 sky130_fd_sc_hd__o2bb2ai_2 _08689_ (.A1_N(_02174_),
    .A2_N(_02175_),
    .B1(_00066_),
    .B2(_00396_),
    .Y(_02682_));
 sky130_fd_sc_hd__o21ai_1 _08690_ (.A1(_00066_),
    .A2(_02176_),
    .B1(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__a31oi_1 _08691_ (.A1(_02655_),
    .A2(net60),
    .A3(net30),
    .B1(_02653_),
    .Y(_02685_));
 sky130_fd_sc_hd__a31o_1 _08692_ (.A1(_02655_),
    .A2(net60),
    .A3(net30),
    .B1(_02653_),
    .X(_02686_));
 sky130_fd_sc_hd__o221ai_4 _08693_ (.A1(_00066_),
    .A2(_02176_),
    .B1(_02653_),
    .B2(_02658_),
    .C1(_02682_),
    .Y(_02687_));
 sky130_fd_sc_hd__nand2_2 _08694_ (.A(_02683_),
    .B(_02685_),
    .Y(_02688_));
 sky130_fd_sc_hd__and3_1 _08695_ (.A(_02681_),
    .B(_02687_),
    .C(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__nand3_4 _08696_ (.A(_02681_),
    .B(_02687_),
    .C(_02688_),
    .Y(_02690_));
 sky130_fd_sc_hd__a21oi_1 _08697_ (.A1(_02687_),
    .A2(_02688_),
    .B1(_02681_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21o_1 _08698_ (.A1(_02687_),
    .A2(_02688_),
    .B1(_02681_),
    .X(_02692_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_02690_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__nand3_2 _08700_ (.A(_02672_),
    .B(_02690_),
    .C(_02692_),
    .Y(_02694_));
 sky130_fd_sc_hd__o21ai_2 _08701_ (.A1(_02671_),
    .A2(_02693_),
    .B1(_02670_),
    .Y(_02696_));
 sky130_fd_sc_hd__o2111ai_4 _08702_ (.A1(_02163_),
    .A2(_02168_),
    .B1(_02194_),
    .C1(_02195_),
    .D1(_02166_),
    .Y(_02697_));
 sky130_fd_sc_hd__o21ai_2 _08703_ (.A1(_02165_),
    .A2(_02169_),
    .B1(_02196_),
    .Y(_02698_));
 sky130_fd_sc_hd__o21ai_2 _08704_ (.A1(_02165_),
    .A2(_02169_),
    .B1(_02197_),
    .Y(_02699_));
 sky130_fd_sc_hd__o2111ai_4 _08705_ (.A1(_02163_),
    .A2(_02168_),
    .B1(_02192_),
    .C1(_02193_),
    .D1(_02166_),
    .Y(_02700_));
 sky130_fd_sc_hd__o2111a_1 _08706_ (.A1(_02665_),
    .A2(_02669_),
    .B1(_02694_),
    .C1(_02697_),
    .D1(_02698_),
    .X(_02701_));
 sky130_fd_sc_hd__o2111ai_4 _08707_ (.A1(_02665_),
    .A2(_02669_),
    .B1(_02694_),
    .C1(_02697_),
    .D1(_02698_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand3_4 _08708_ (.A(_02696_),
    .B(_02699_),
    .C(_02700_),
    .Y(_02703_));
 sky130_fd_sc_hd__o22ai_4 _08709_ (.A1(_00055_),
    .A2(_00407_),
    .B1(_02309_),
    .B2(_02311_),
    .Y(_02704_));
 sky130_fd_sc_hd__a22oi_2 _08710_ (.A1(net26),
    .A2(net64),
    .B1(net34),
    .B2(net23),
    .Y(_02705_));
 sky130_fd_sc_hd__a22o_1 _08711_ (.A1(net26),
    .A2(net64),
    .B1(net34),
    .B2(net23),
    .X(_02707_));
 sky130_fd_sc_hd__and4_1 _08712_ (.A(net26),
    .B(net23),
    .C(net64),
    .D(net34),
    .X(_02708_));
 sky130_fd_sc_hd__nand4_4 _08713_ (.A(net26),
    .B(net23),
    .C(net64),
    .D(net34),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(net12),
    .B(net35),
    .Y(_02710_));
 sky130_fd_sc_hd__o21ai_4 _08715_ (.A1(_02710_),
    .A2(_02705_),
    .B1(_02709_),
    .Y(_02711_));
 sky130_fd_sc_hd__and3_1 _08716_ (.A(_02313_),
    .B(_02704_),
    .C(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__nand3_4 _08717_ (.A(_02313_),
    .B(_02704_),
    .C(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hd__and4_2 _08718_ (.A(net12),
    .B(net1),
    .C(net37),
    .D(net36),
    .X(_02714_));
 sky130_fd_sc_hd__nand4_1 _08719_ (.A(net12),
    .B(net1),
    .C(net37),
    .D(net36),
    .Y(_02715_));
 sky130_fd_sc_hd__o2bb2a_1 _08720_ (.A1_N(net1),
    .A2_N(net37),
    .B1(_00429_),
    .B2(_00022_),
    .X(_02716_));
 sky130_fd_sc_hd__nor2_1 _08721_ (.A(_02714_),
    .B(_02716_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21oi_1 _08722_ (.A1(_02313_),
    .A2(_02704_),
    .B1(_02711_),
    .Y(_02719_));
 sky130_fd_sc_hd__a21o_1 _08723_ (.A1(_02313_),
    .A2(_02704_),
    .B1(_02711_),
    .X(_02720_));
 sky130_fd_sc_hd__nand3_4 _08724_ (.A(_02713_),
    .B(_02720_),
    .C(_02718_),
    .Y(_02721_));
 sky130_fd_sc_hd__a21o_1 _08725_ (.A1(_02720_),
    .A2(_02718_),
    .B1(_02712_),
    .X(_02722_));
 sky130_fd_sc_hd__o211ai_2 _08726_ (.A1(_02324_),
    .A2(_02325_),
    .B1(_02318_),
    .C1(_02319_),
    .Y(_02723_));
 sky130_fd_sc_hd__o2bb2ai_2 _08727_ (.A1_N(_02318_),
    .A2_N(_02319_),
    .B1(_02326_),
    .B2(_02327_),
    .Y(_02724_));
 sky130_fd_sc_hd__o2bb2ai_1 _08728_ (.A1_N(_02318_),
    .A2_N(_02319_),
    .B1(_02324_),
    .B2(_02325_),
    .Y(_02725_));
 sky130_fd_sc_hd__o211ai_2 _08729_ (.A1(_02326_),
    .A2(_02327_),
    .B1(_02318_),
    .C1(_02319_),
    .Y(_02726_));
 sky130_fd_sc_hd__a32o_1 _08730_ (.A1(_02177_),
    .A2(_02682_),
    .A3(_02686_),
    .B1(_02688_),
    .B2(_02681_),
    .X(_02727_));
 sky130_fd_sc_hd__a21oi_2 _08731_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__a21o_1 _08732_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02727_),
    .X(_02730_));
 sky130_fd_sc_hd__a22oi_4 _08733_ (.A1(_02687_),
    .A2(_02690_),
    .B1(_02723_),
    .B2(_02724_),
    .Y(_02731_));
 sky130_fd_sc_hd__a22o_1 _08734_ (.A1(_02687_),
    .A2(_02690_),
    .B1(_02723_),
    .B2(_02724_),
    .X(_02732_));
 sky130_fd_sc_hd__a211oi_4 _08735_ (.A1(_02713_),
    .A2(_02721_),
    .B1(_02729_),
    .C1(_02731_),
    .Y(_02733_));
 sky130_fd_sc_hd__nand3_2 _08736_ (.A(_02722_),
    .B(_02730_),
    .C(_02732_),
    .Y(_02734_));
 sky130_fd_sc_hd__o211a_1 _08737_ (.A1(_02729_),
    .A2(_02731_),
    .B1(_02713_),
    .C1(_02721_),
    .X(_02735_));
 sky130_fd_sc_hd__o211ai_2 _08738_ (.A1(_02729_),
    .A2(_02731_),
    .B1(_02713_),
    .C1(_02721_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_1 _08739_ (.A(_02734_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__a32oi_1 _08740_ (.A1(_02696_),
    .A2(_02699_),
    .A3(_02700_),
    .B1(_02734_),
    .B2(_02736_),
    .Y(_02738_));
 sky130_fd_sc_hd__a32o_1 _08741_ (.A1(_02696_),
    .A2(_02699_),
    .A3(_02700_),
    .B1(_02734_),
    .B2(_02736_),
    .X(_02740_));
 sky130_fd_sc_hd__o211ai_2 _08742_ (.A1(_02261_),
    .A2(_02267_),
    .B1(_02270_),
    .C1(_02333_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _08743_ (.A(_02269_),
    .B(_02270_),
    .Y(_02742_));
 sky130_fd_sc_hd__o2bb2ai_2 _08744_ (.A1_N(_02269_),
    .A2_N(_02270_),
    .B1(_02330_),
    .B2(_02331_),
    .Y(_02743_));
 sky130_fd_sc_hd__o221ai_4 _08745_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_02261_),
    .B2(_02267_),
    .C1(_02270_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand2_1 _08746_ (.A(_02742_),
    .B(_02333_),
    .Y(_02745_));
 sky130_fd_sc_hd__a2bb2oi_1 _08747_ (.A1_N(_02701_),
    .A2_N(_02738_),
    .B1(_02741_),
    .B2(_02743_),
    .Y(_02746_));
 sky130_fd_sc_hd__o2111ai_4 _08748_ (.A1(_02737_),
    .A2(_02701_),
    .B1(_02703_),
    .C1(_02744_),
    .D1(_02745_),
    .Y(_02747_));
 sky130_fd_sc_hd__o2111a_1 _08749_ (.A1(_02268_),
    .A2(_02334_),
    .B1(_02702_),
    .C1(_02740_),
    .D1(_02743_),
    .X(_02748_));
 sky130_fd_sc_hd__o2111ai_4 _08750_ (.A1(_02268_),
    .A2(_02334_),
    .B1(_02702_),
    .C1(_02740_),
    .D1(_02743_),
    .Y(_02749_));
 sky130_fd_sc_hd__a21oi_2 _08751_ (.A1(_02722_),
    .A2(_02730_),
    .B1(_02731_),
    .Y(_02751_));
 sky130_fd_sc_hd__a211o_1 _08752_ (.A1(net1),
    .A2(net39),
    .B1(_02320_),
    .C1(_02324_),
    .X(_02752_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(_02441_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__o211a_1 _08754_ (.A1(_02731_),
    .A2(_02733_),
    .B1(_02752_),
    .C1(_02441_),
    .X(_02754_));
 sky130_fd_sc_hd__o21bai_2 _08755_ (.A1(_02731_),
    .A2(_02733_),
    .B1_N(_02753_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_02751_),
    .B(_02753_),
    .Y(_02756_));
 sky130_fd_sc_hd__and2_1 _08757_ (.A(_02755_),
    .B(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__nand2_1 _08758_ (.A(_02755_),
    .B(_02756_),
    .Y(_02758_));
 sky130_fd_sc_hd__a41o_1 _08759_ (.A1(_02702_),
    .A2(_02740_),
    .A3(_02741_),
    .A4(_02743_),
    .B1(_02757_),
    .X(_02759_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_02747_),
    .B(_02757_),
    .Y(_02760_));
 sky130_fd_sc_hd__a22oi_2 _08761_ (.A1(_02452_),
    .A2(_02454_),
    .B1(_02457_),
    .B2(_02437_),
    .Y(_02762_));
 sky130_fd_sc_hd__a22o_1 _08762_ (.A1(_02452_),
    .A2(_02454_),
    .B1(_02457_),
    .B2(_02437_),
    .X(_02763_));
 sky130_fd_sc_hd__a221oi_2 _08763_ (.A1(_02458_),
    .A2(_02437_),
    .B1(_02760_),
    .B2(_02749_),
    .C1(_02762_),
    .Y(_02764_));
 sky130_fd_sc_hd__o2111ai_2 _08764_ (.A1(_02436_),
    .A2(_02459_),
    .B1(_02747_),
    .C1(_02759_),
    .D1(_02763_),
    .Y(_02765_));
 sky130_fd_sc_hd__a22oi_2 _08765_ (.A1(_02747_),
    .A2(_02759_),
    .B1(_02763_),
    .B2(_02461_),
    .Y(_02766_));
 sky130_fd_sc_hd__o2bb2ai_1 _08766_ (.A1_N(_02747_),
    .A2_N(_02759_),
    .B1(_02762_),
    .B2(_02460_),
    .Y(_02767_));
 sky130_fd_sc_hd__o21ai_1 _08767_ (.A1(_02755_),
    .A2(_02766_),
    .B1(_02765_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand3_1 _08768_ (.A(_02565_),
    .B(_02638_),
    .C(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__a22oi_4 _08769_ (.A1(net32),
    .A2(net44),
    .B1(net33),
    .B2(net2),
    .Y(_02770_));
 sky130_fd_sc_hd__a22o_1 _08770_ (.A1(net32),
    .A2(net44),
    .B1(net33),
    .B2(net2),
    .X(_02771_));
 sky130_fd_sc_hd__and4_1 _08771_ (.A(net32),
    .B(net2),
    .C(net44),
    .D(net33),
    .X(_02773_));
 sky130_fd_sc_hd__nand4_4 _08772_ (.A(net32),
    .B(net2),
    .C(net44),
    .D(net33),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(net31),
    .B(net55),
    .Y(_02775_));
 sky130_fd_sc_hd__o21ai_2 _08774_ (.A1(_02775_),
    .A2(_02770_),
    .B1(_02774_),
    .Y(_02776_));
 sky130_fd_sc_hd__o21a_1 _08775_ (.A1(_02775_),
    .A2(_02770_),
    .B1(_02774_),
    .X(_02777_));
 sky130_fd_sc_hd__o211ai_1 _08776_ (.A1(_00110_),
    .A2(_00341_),
    .B1(_02642_),
    .C1(_02644_),
    .Y(_02778_));
 sky130_fd_sc_hd__o21bai_1 _08777_ (.A1(_02641_),
    .A2(_02643_),
    .B1_N(_02645_),
    .Y(_02779_));
 sky130_fd_sc_hd__o22a_1 _08778_ (.A1(_00110_),
    .A2(_00341_),
    .B1(_02641_),
    .B2(_02643_),
    .X(_02780_));
 sky130_fd_sc_hd__o22ai_2 _08779_ (.A1(_00110_),
    .A2(_00341_),
    .B1(_02641_),
    .B2(_02643_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand4_2 _08780_ (.A(_02642_),
    .B(_02644_),
    .C(net32),
    .D(net55),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_1 _08781_ (.A(_02776_),
    .B(_02782_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand3_2 _08782_ (.A(_02781_),
    .B(_02782_),
    .C(_02776_),
    .Y(_02785_));
 sky130_fd_sc_hd__a21oi_2 _08783_ (.A1(_02781_),
    .A2(_02782_),
    .B1(_02776_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand3_2 _08784_ (.A(_02777_),
    .B(_02778_),
    .C(_02779_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_1 _08785_ (.A(net29),
    .B(net60),
    .Y(_02788_));
 sky130_fd_sc_hd__and4_1 _08786_ (.A(net30),
    .B(net31),
    .C(net58),
    .D(net59),
    .X(_02789_));
 sky130_fd_sc_hd__nand4_2 _08787_ (.A(net30),
    .B(net31),
    .C(net58),
    .D(net59),
    .Y(_02790_));
 sky130_fd_sc_hd__a22oi_2 _08788_ (.A1(net31),
    .A2(net58),
    .B1(net59),
    .B2(net30),
    .Y(_02791_));
 sky130_fd_sc_hd__a22o_1 _08789_ (.A1(net31),
    .A2(net58),
    .B1(net59),
    .B2(net30),
    .X(_02792_));
 sky130_fd_sc_hd__o22a_1 _08790_ (.A1(_00099_),
    .A2(_00352_),
    .B1(_02789_),
    .B2(_02791_),
    .X(_02793_));
 sky130_fd_sc_hd__o22ai_2 _08791_ (.A1(_00099_),
    .A2(_00352_),
    .B1(_02789_),
    .B2(_02791_),
    .Y(_02795_));
 sky130_fd_sc_hd__and4_1 _08792_ (.A(_02792_),
    .B(net60),
    .C(net29),
    .D(_02790_),
    .X(_02796_));
 sky130_fd_sc_hd__nand4_2 _08793_ (.A(_02792_),
    .B(net60),
    .C(net29),
    .D(_02790_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_02795_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand4_4 _08795_ (.A(_02785_),
    .B(_02787_),
    .C(_02795_),
    .D(_02797_),
    .Y(_02799_));
 sky130_fd_sc_hd__o22a_1 _08796_ (.A1(_02784_),
    .A2(_02780_),
    .B1(_02798_),
    .B2(_02786_),
    .X(_02800_));
 sky130_fd_sc_hd__o22ai_4 _08797_ (.A1(_02784_),
    .A2(_02780_),
    .B1(_02798_),
    .B2(_02786_),
    .Y(_02801_));
 sky130_fd_sc_hd__o22ai_4 _08798_ (.A1(_02656_),
    .A2(_02658_),
    .B1(_02660_),
    .B2(_02652_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _08799_ (.A(_02664_),
    .B(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__a21oi_2 _08800_ (.A1(_02664_),
    .A2(_02802_),
    .B1(_02801_),
    .Y(_02804_));
 sky130_fd_sc_hd__a21o_1 _08801_ (.A1(_02664_),
    .A2(_02802_),
    .B1(_02801_),
    .X(_02806_));
 sky130_fd_sc_hd__nand2_1 _08802_ (.A(_02801_),
    .B(_02802_),
    .Y(_02807_));
 sky130_fd_sc_hd__and3_1 _08803_ (.A(_02664_),
    .B(_02801_),
    .C(_02802_),
    .X(_02808_));
 sky130_fd_sc_hd__nand2_1 _08804_ (.A(_02788_),
    .B(_02790_),
    .Y(_02809_));
 sky130_fd_sc_hd__o211ai_2 _08805_ (.A1(_00077_),
    .A2(_00396_),
    .B1(_02678_),
    .C1(_02679_),
    .Y(_02810_));
 sky130_fd_sc_hd__and4_1 _08806_ (.A(_02680_),
    .B(_02792_),
    .C(_02809_),
    .D(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__nand4_1 _08807_ (.A(_02680_),
    .B(_02792_),
    .C(_02809_),
    .D(_02810_),
    .Y(_02812_));
 sky130_fd_sc_hd__a22o_1 _08808_ (.A1(_02792_),
    .A2(_02809_),
    .B1(_02810_),
    .B2(_02680_),
    .X(_02813_));
 sky130_fd_sc_hd__o22a_1 _08809_ (.A1(_00077_),
    .A2(_00374_),
    .B1(_00385_),
    .B2(_00066_),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_1 _08810_ (.A1(net27),
    .A2(net62),
    .B1(net61),
    .B2(net28),
    .X(_02815_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(net27),
    .B(net61),
    .Y(_02817_));
 sky130_fd_sc_hd__and4_1 _08812_ (.A(net28),
    .B(net27),
    .C(net62),
    .D(net61),
    .X(_02818_));
 sky130_fd_sc_hd__nand4_1 _08813_ (.A(net28),
    .B(net27),
    .C(net62),
    .D(net61),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(net26),
    .B(net63),
    .Y(_02820_));
 sky130_fd_sc_hd__and3_1 _08815_ (.A(_02815_),
    .B(net63),
    .C(net26),
    .X(_02821_));
 sky130_fd_sc_hd__a31o_1 _08816_ (.A1(_02815_),
    .A2(net63),
    .A3(net26),
    .B1(_02818_),
    .X(_02822_));
 sky130_fd_sc_hd__o211a_2 _08817_ (.A1(_02818_),
    .A2(_02821_),
    .B1(_02812_),
    .C1(_02813_),
    .X(_02823_));
 sky130_fd_sc_hd__a21oi_2 _08818_ (.A1(_02812_),
    .A2(_02813_),
    .B1(_02822_),
    .Y(_02824_));
 sky130_fd_sc_hd__nor2_1 _08819_ (.A(_02823_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__o22a_1 _08820_ (.A1(_02823_),
    .A2(_02824_),
    .B1(_02800_),
    .B2(_02803_),
    .X(_02826_));
 sky130_fd_sc_hd__a211oi_1 _08821_ (.A1(_02803_),
    .A2(_02800_),
    .B1(_02824_),
    .C1(_02823_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand4_2 _08822_ (.A(_02670_),
    .B(_02672_),
    .C(_02690_),
    .D(_02692_),
    .Y(_02829_));
 sky130_fd_sc_hd__o2bb2ai_2 _08823_ (.A1_N(_02670_),
    .A2_N(_02672_),
    .B1(_02689_),
    .B2(_02691_),
    .Y(_02830_));
 sky130_fd_sc_hd__o211ai_1 _08824_ (.A1(_02689_),
    .A2(_02691_),
    .B1(_02670_),
    .C1(_02672_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21o_1 _08825_ (.A1(_02670_),
    .A2(_02672_),
    .B1(_02693_),
    .X(_02832_));
 sky130_fd_sc_hd__o211a_1 _08826_ (.A1(_02808_),
    .A2(_02828_),
    .B1(_02829_),
    .C1(_02830_),
    .X(_02833_));
 sky130_fd_sc_hd__o211ai_2 _08827_ (.A1(_02808_),
    .A2(_02828_),
    .B1(_02829_),
    .C1(_02830_),
    .Y(_02834_));
 sky130_fd_sc_hd__and4_2 _08828_ (.A(net12),
    .B(net23),
    .C(net64),
    .D(net34),
    .X(_02835_));
 sky130_fd_sc_hd__nand4_2 _08829_ (.A(net12),
    .B(net23),
    .C(net64),
    .D(net34),
    .Y(_02836_));
 sky130_fd_sc_hd__a22o_1 _08830_ (.A1(net23),
    .A2(net64),
    .B1(net34),
    .B2(net12),
    .X(_02837_));
 sky130_fd_sc_hd__nand4_4 _08831_ (.A(_02837_),
    .B(net35),
    .C(net1),
    .D(_02836_),
    .Y(_02839_));
 sky130_fd_sc_hd__a31o_1 _08832_ (.A1(_02837_),
    .A2(net35),
    .A3(net1),
    .B1(_02835_),
    .X(_02840_));
 sky130_fd_sc_hd__o211ai_1 _08833_ (.A1(_00022_),
    .A2(_00407_),
    .B1(_02707_),
    .C1(_02709_),
    .Y(_02841_));
 sky130_fd_sc_hd__o21bai_1 _08834_ (.A1(_02705_),
    .A2(_02708_),
    .B1_N(_02710_),
    .Y(_02842_));
 sky130_fd_sc_hd__a22o_1 _08835_ (.A1(net12),
    .A2(net35),
    .B1(_02707_),
    .B2(_02709_),
    .X(_02843_));
 sky130_fd_sc_hd__nand4_2 _08836_ (.A(_02707_),
    .B(_02709_),
    .C(net12),
    .D(net35),
    .Y(_02844_));
 sky130_fd_sc_hd__nand3_2 _08837_ (.A(_02839_),
    .B(_02841_),
    .C(_02842_),
    .Y(_02845_));
 sky130_fd_sc_hd__nor2_1 _08838_ (.A(_02835_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__and3_1 _08839_ (.A(_02840_),
    .B(_02843_),
    .C(_02844_),
    .X(_02847_));
 sky130_fd_sc_hd__nand3_2 _08840_ (.A(_02840_),
    .B(_02843_),
    .C(_02844_),
    .Y(_02848_));
 sky130_fd_sc_hd__o21a_1 _08841_ (.A1(_00033_),
    .A2(_00429_),
    .B1(_02848_),
    .X(_02850_));
 sky130_fd_sc_hd__o211a_1 _08842_ (.A1(_02835_),
    .A2(_02845_),
    .B1(net1),
    .C1(net36),
    .X(_02851_));
 sky130_fd_sc_hd__a31o_1 _08843_ (.A1(_02840_),
    .A2(_02843_),
    .A3(_02844_),
    .B1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a21o_1 _08844_ (.A1(_02813_),
    .A2(_02822_),
    .B1(_02811_),
    .X(_02853_));
 sky130_fd_sc_hd__o22ai_2 _08845_ (.A1(_02714_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02712_),
    .Y(_02854_));
 sky130_fd_sc_hd__o211a_1 _08846_ (.A1(_02811_),
    .A2(_02823_),
    .B1(_02854_),
    .C1(_02721_),
    .X(_02855_));
 sky130_fd_sc_hd__o211ai_1 _08847_ (.A1(_02811_),
    .A2(_02823_),
    .B1(_02854_),
    .C1(_02721_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21oi_1 _08848_ (.A1(_02721_),
    .A2(_02854_),
    .B1(_02853_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21o_1 _08849_ (.A1(_02721_),
    .A2(_02854_),
    .B1(_02853_),
    .X(_02858_));
 sky130_fd_sc_hd__and3_1 _08850_ (.A(_02858_),
    .B(_02852_),
    .C(_02856_),
    .X(_02859_));
 sky130_fd_sc_hd__o211ai_2 _08851_ (.A1(_02847_),
    .A2(_02851_),
    .B1(_02856_),
    .C1(_02858_),
    .Y(_02861_));
 sky130_fd_sc_hd__o22a_1 _08852_ (.A1(_02846_),
    .A2(_02850_),
    .B1(_02855_),
    .B2(_02857_),
    .X(_02862_));
 sky130_fd_sc_hd__o22ai_2 _08853_ (.A1(_02846_),
    .A2(_02850_),
    .B1(_02855_),
    .B2(_02857_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_02861_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__a2bb2oi_2 _08855_ (.A1_N(_02804_),
    .A2_N(_02826_),
    .B1(_02829_),
    .B2(_02830_),
    .Y(_02865_));
 sky130_fd_sc_hd__o211ai_1 _08856_ (.A1(_02804_),
    .A2(_02826_),
    .B1(_02831_),
    .C1(_02832_),
    .Y(_02866_));
 sky130_fd_sc_hd__nand4_2 _08857_ (.A(_02834_),
    .B(_02861_),
    .C(_02863_),
    .D(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__o21a_1 _08858_ (.A1(_02864_),
    .A2(_02865_),
    .B1(_02834_),
    .X(_02868_));
 sky130_fd_sc_hd__o21ai_1 _08859_ (.A1(_02864_),
    .A2(_02865_),
    .B1(_02834_),
    .Y(_02869_));
 sky130_fd_sc_hd__o211ai_2 _08860_ (.A1(_02733_),
    .A2(_02735_),
    .B1(_02702_),
    .C1(_02703_),
    .Y(_02870_));
 sky130_fd_sc_hd__a21o_1 _08861_ (.A1(_02702_),
    .A2(_02703_),
    .B1(_02737_),
    .X(_02872_));
 sky130_fd_sc_hd__nand4_1 _08862_ (.A(_02702_),
    .B(_02703_),
    .C(_02734_),
    .D(_02736_),
    .Y(_02873_));
 sky130_fd_sc_hd__o2bb2ai_1 _08863_ (.A1_N(_02702_),
    .A2_N(_02703_),
    .B1(_02733_),
    .B2(_02735_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand3_1 _08864_ (.A(_02872_),
    .B(_02868_),
    .C(_02870_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand3_2 _08865_ (.A(_02869_),
    .B(_02873_),
    .C(_02874_),
    .Y(_02876_));
 sky130_fd_sc_hd__a21o_2 _08866_ (.A1(_02858_),
    .A2(_02852_),
    .B1(_02855_),
    .X(_02877_));
 sky130_fd_sc_hd__inv_2 _08867_ (.A(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__xor2_1 _08868_ (.A(_02714_),
    .B(_02877_),
    .X(_02879_));
 sky130_fd_sc_hd__xor2_1 _08869_ (.A(_02715_),
    .B(_02877_),
    .X(_02880_));
 sky130_fd_sc_hd__a32oi_2 _08870_ (.A1(_02868_),
    .A2(_02870_),
    .A3(_02872_),
    .B1(_02876_),
    .B2(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__a32o_1 _08871_ (.A1(_02868_),
    .A2(_02870_),
    .A3(_02872_),
    .B1(_02876_),
    .B2(_02880_),
    .X(_02883_));
 sky130_fd_sc_hd__o21bai_1 _08872_ (.A1(_02746_),
    .A2(_02748_),
    .B1_N(_02758_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand3_1 _08873_ (.A(_02747_),
    .B(_02749_),
    .C(_02758_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand4_1 _08874_ (.A(_02747_),
    .B(_02749_),
    .C(_02755_),
    .D(_02756_),
    .Y(_02886_));
 sky130_fd_sc_hd__o21ai_1 _08875_ (.A1(_02746_),
    .A2(_02748_),
    .B1(_02758_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand3_1 _08876_ (.A(_02887_),
    .B(_02881_),
    .C(_02886_),
    .Y(_02888_));
 sky130_fd_sc_hd__o22ai_1 _08877_ (.A1(_02751_),
    .A2(_02753_),
    .B1(_02764_),
    .B2(_02766_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand3_1 _08878_ (.A(_02767_),
    .B(_02754_),
    .C(_02765_),
    .Y(_02890_));
 sky130_fd_sc_hd__o21bai_1 _08879_ (.A1(_02764_),
    .A2(_02766_),
    .B1_N(_02755_),
    .Y(_02891_));
 sky130_fd_sc_hd__o211ai_1 _08880_ (.A1(_02751_),
    .A2(_02753_),
    .B1(_02765_),
    .C1(_02767_),
    .Y(_02892_));
 sky130_fd_sc_hd__a32o_1 _08881_ (.A1(_02887_),
    .A2(_02881_),
    .A3(_02886_),
    .B1(_02877_),
    .B2(_02714_),
    .X(_02894_));
 sky130_fd_sc_hd__nand3_1 _08882_ (.A(_02883_),
    .B(_02884_),
    .C(_02885_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand4_1 _08883_ (.A(_02889_),
    .B(_02890_),
    .C(_02894_),
    .D(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__a22oi_4 _08884_ (.A1(net29),
    .A2(net58),
    .B1(net59),
    .B2(net28),
    .Y(_02897_));
 sky130_fd_sc_hd__a22o_1 _08885_ (.A1(net29),
    .A2(net58),
    .B1(net59),
    .B2(net28),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(net27),
    .B(net60),
    .Y(_02899_));
 sky130_fd_sc_hd__and4_1 _08887_ (.A(net28),
    .B(net29),
    .C(net58),
    .D(net59),
    .X(_02900_));
 sky130_fd_sc_hd__nand4_4 _08888_ (.A(net28),
    .B(net29),
    .C(net58),
    .D(net59),
    .Y(_02901_));
 sky130_fd_sc_hd__o21ai_4 _08889_ (.A1(_02899_),
    .A2(_02897_),
    .B1(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(net26),
    .B(net62),
    .Y(_02903_));
 sky130_fd_sc_hd__and4_1 _08891_ (.A(net26),
    .B(net27),
    .C(net62),
    .D(net61),
    .X(_02905_));
 sky130_fd_sc_hd__nand4_1 _08892_ (.A(net26),
    .B(net27),
    .C(net62),
    .D(net61),
    .Y(_02906_));
 sky130_fd_sc_hd__a22o_1 _08893_ (.A1(net26),
    .A2(net62),
    .B1(net61),
    .B2(net27),
    .X(_02907_));
 sky130_fd_sc_hd__nand3_1 _08894_ (.A(_02903_),
    .B(net61),
    .C(net27),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _08895_ (.A(_02817_),
    .B(net62),
    .C(net26),
    .Y(_02909_));
 sky130_fd_sc_hd__and4_1 _08896_ (.A(_02907_),
    .B(net63),
    .C(net23),
    .D(_02906_),
    .X(_02910_));
 sky130_fd_sc_hd__nand4_2 _08897_ (.A(_02907_),
    .B(net63),
    .C(net23),
    .D(_02906_),
    .Y(_02911_));
 sky130_fd_sc_hd__o211ai_4 _08898_ (.A1(_00055_),
    .A2(_00396_),
    .B1(_02908_),
    .C1(_02909_),
    .Y(_02912_));
 sky130_fd_sc_hd__and3_2 _08899_ (.A(_02912_),
    .B(_02902_),
    .C(_02911_),
    .X(_02913_));
 sky130_fd_sc_hd__nand3_1 _08900_ (.A(_02902_),
    .B(_02911_),
    .C(_02912_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand4_4 _08901_ (.A(net26),
    .B(net23),
    .C(net62),
    .D(net61),
    .Y(_02916_));
 sky130_fd_sc_hd__a22o_1 _08902_ (.A1(net23),
    .A2(net62),
    .B1(net61),
    .B2(net26),
    .X(_02917_));
 sky130_fd_sc_hd__nand4_4 _08903_ (.A(_02917_),
    .B(net63),
    .C(net12),
    .D(_02916_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(_02916_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21oi_2 _08905_ (.A1(_02911_),
    .A2(_02912_),
    .B1(_02902_),
    .Y(_02920_));
 sky130_fd_sc_hd__a21o_1 _08906_ (.A1(_02911_),
    .A2(_02912_),
    .B1(_02902_),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(_02919_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__a211o_2 _08908_ (.A1(_02916_),
    .A2(_02918_),
    .B1(_02920_),
    .C1(_02913_),
    .X(_02923_));
 sky130_fd_sc_hd__a21oi_2 _08909_ (.A1(_02919_),
    .A2(_02921_),
    .B1(_02913_),
    .Y(_02924_));
 sky130_fd_sc_hd__and4_1 _08910_ (.A(net12),
    .B(net1),
    .C(net64),
    .D(net34),
    .X(_02925_));
 sky130_fd_sc_hd__nand4_2 _08911_ (.A(net12),
    .B(net1),
    .C(net64),
    .D(net34),
    .Y(_02927_));
 sky130_fd_sc_hd__a22o_1 _08912_ (.A1(net1),
    .A2(net35),
    .B1(_02836_),
    .B2(_02837_),
    .X(_02928_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_02839_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__and3_1 _08914_ (.A(_02839_),
    .B(_02928_),
    .C(_02925_),
    .X(_02930_));
 sky130_fd_sc_hd__nand3_1 _08915_ (.A(_02839_),
    .B(_02928_),
    .C(_02925_),
    .Y(_02931_));
 sky130_fd_sc_hd__a21o_1 _08916_ (.A1(_02839_),
    .A2(_02928_),
    .B1(_02925_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_2 _08917_ (.A(_02931_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__a21oi_1 _08918_ (.A1(_02914_),
    .A2(_02923_),
    .B1(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__a21o_1 _08919_ (.A1(_02914_),
    .A2(_02923_),
    .B1(_02933_),
    .X(_02935_));
 sky130_fd_sc_hd__a31o_1 _08920_ (.A1(_02907_),
    .A2(net63),
    .A3(net23),
    .B1(_02905_),
    .X(_02936_));
 sky130_fd_sc_hd__a22oi_4 _08921_ (.A1(net30),
    .A2(net58),
    .B1(net59),
    .B2(net29),
    .Y(_02938_));
 sky130_fd_sc_hd__a22o_1 _08922_ (.A1(net30),
    .A2(net58),
    .B1(net59),
    .B2(net29),
    .X(_02939_));
 sky130_fd_sc_hd__and4_2 _08923_ (.A(net30),
    .B(net29),
    .C(net58),
    .D(net59),
    .X(_02940_));
 sky130_fd_sc_hd__a31o_1 _08924_ (.A1(_02939_),
    .A2(net60),
    .A3(net28),
    .B1(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__a31oi_1 _08925_ (.A1(_02939_),
    .A2(net60),
    .A3(net28),
    .B1(_02940_),
    .Y(_02942_));
 sky130_fd_sc_hd__o221ai_2 _08926_ (.A1(_00044_),
    .A2(_00396_),
    .B1(_02675_),
    .B2(_02817_),
    .C1(_02815_),
    .Y(_02943_));
 sky130_fd_sc_hd__a21o_1 _08927_ (.A1(_02815_),
    .A2(_02819_),
    .B1(_02820_),
    .X(_02944_));
 sky130_fd_sc_hd__a41o_1 _08928_ (.A1(net28),
    .A2(net27),
    .A3(net62),
    .A4(net61),
    .B1(_02820_),
    .X(_02945_));
 sky130_fd_sc_hd__and4_1 _08929_ (.A(_02815_),
    .B(_02819_),
    .C(net26),
    .D(net63),
    .X(_02946_));
 sky130_fd_sc_hd__a22o_1 _08930_ (.A1(net26),
    .A2(net63),
    .B1(_02815_),
    .B2(_02819_),
    .X(_02947_));
 sky130_fd_sc_hd__nand2_1 _08931_ (.A(_02941_),
    .B(_02947_),
    .Y(_02949_));
 sky130_fd_sc_hd__o211ai_4 _08932_ (.A1(_02945_),
    .A2(_02814_),
    .B1(_02947_),
    .C1(_02941_),
    .Y(_02950_));
 sky130_fd_sc_hd__nand3_2 _08933_ (.A(_02942_),
    .B(_02943_),
    .C(_02944_),
    .Y(_02951_));
 sky130_fd_sc_hd__o21a_1 _08934_ (.A1(_02905_),
    .A2(_02910_),
    .B1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__o221a_2 _08935_ (.A1(_02905_),
    .A2(_02910_),
    .B1(_02946_),
    .B2(_02949_),
    .C1(_02951_),
    .X(_02953_));
 sky130_fd_sc_hd__a21oi_4 _08936_ (.A1(_02950_),
    .A2(_02951_),
    .B1(_02936_),
    .Y(_02954_));
 sky130_fd_sc_hd__a21oi_2 _08937_ (.A1(_02952_),
    .A2(_02950_),
    .B1(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__a22oi_4 _08938_ (.A1(net31),
    .A2(net44),
    .B1(net33),
    .B2(net32),
    .Y(_02956_));
 sky130_fd_sc_hd__a22o_1 _08939_ (.A1(net31),
    .A2(net44),
    .B1(net33),
    .B2(net32),
    .X(_02957_));
 sky130_fd_sc_hd__and4_1 _08940_ (.A(net32),
    .B(net31),
    .C(net44),
    .D(net33),
    .X(_02958_));
 sky130_fd_sc_hd__nand4_4 _08941_ (.A(net32),
    .B(net31),
    .C(net44),
    .D(net33),
    .Y(_02960_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(net30),
    .B(net55),
    .Y(_02961_));
 sky130_fd_sc_hd__o21ai_2 _08943_ (.A1(_02961_),
    .A2(_02956_),
    .B1(_02960_),
    .Y(_02962_));
 sky130_fd_sc_hd__o21a_2 _08944_ (.A1(_02961_),
    .A2(_02956_),
    .B1(_02960_),
    .X(_02963_));
 sky130_fd_sc_hd__o211ai_4 _08945_ (.A1(_00121_),
    .A2(_00341_),
    .B1(_02771_),
    .C1(_02774_),
    .Y(_02964_));
 sky130_fd_sc_hd__o21bai_4 _08946_ (.A1(_02770_),
    .A2(_02773_),
    .B1_N(_02775_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand4_2 _08947_ (.A(_02771_),
    .B(_02774_),
    .C(net31),
    .D(net55),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_2 _08948_ (.A1(_02770_),
    .A2(_02773_),
    .B1(_02775_),
    .Y(_02967_));
 sky130_fd_sc_hd__nand3_4 _08949_ (.A(_02963_),
    .B(_02964_),
    .C(_02965_),
    .Y(_02968_));
 sky130_fd_sc_hd__and3_2 _08950_ (.A(_02967_),
    .B(_02962_),
    .C(_02966_),
    .X(_02969_));
 sky130_fd_sc_hd__nand3_4 _08951_ (.A(_02967_),
    .B(_02962_),
    .C(_02966_),
    .Y(_02971_));
 sky130_fd_sc_hd__a211oi_2 _08952_ (.A1(net28),
    .A2(net60),
    .B1(_02938_),
    .C1(_02940_),
    .Y(_02972_));
 sky130_fd_sc_hd__a211o_2 _08953_ (.A1(net28),
    .A2(net60),
    .B1(_02938_),
    .C1(_02940_),
    .X(_02973_));
 sky130_fd_sc_hd__o211a_1 _08954_ (.A1(_02938_),
    .A2(_02940_),
    .B1(net28),
    .C1(net60),
    .X(_02974_));
 sky130_fd_sc_hd__o211ai_4 _08955_ (.A1(_02938_),
    .A2(_02940_),
    .B1(net28),
    .C1(net60),
    .Y(_02975_));
 sky130_fd_sc_hd__o22a_1 _08956_ (.A1(_00066_),
    .A2(_00352_),
    .B1(_02938_),
    .B2(_02940_),
    .X(_02976_));
 sky130_fd_sc_hd__and4b_1 _08957_ (.A_N(_02940_),
    .B(net60),
    .C(net28),
    .D(_02939_),
    .X(_02977_));
 sky130_fd_sc_hd__nand3_2 _08958_ (.A(_02971_),
    .B(_02973_),
    .C(_02975_),
    .Y(_02978_));
 sky130_fd_sc_hd__a32oi_4 _08959_ (.A1(_02963_),
    .A2(_02964_),
    .A3(_02965_),
    .B1(_02973_),
    .B2(_02975_),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_1 _08960_ (.A1(_02972_),
    .A2(_02974_),
    .B1(_02968_),
    .Y(_02980_));
 sky130_fd_sc_hd__o2bb2ai_4 _08961_ (.A1_N(_02785_),
    .A2_N(_02787_),
    .B1(_02793_),
    .B2(_02796_),
    .Y(_02982_));
 sky130_fd_sc_hd__o211a_2 _08962_ (.A1(_02969_),
    .A2(_02979_),
    .B1(_02982_),
    .C1(_02799_),
    .X(_02983_));
 sky130_fd_sc_hd__o211ai_4 _08963_ (.A1(_02969_),
    .A2(_02979_),
    .B1(_02982_),
    .C1(_02799_),
    .Y(_02984_));
 sky130_fd_sc_hd__a22oi_4 _08964_ (.A1(_02968_),
    .A2(_02978_),
    .B1(_02982_),
    .B2(_02799_),
    .Y(_02985_));
 sky130_fd_sc_hd__a22o_2 _08965_ (.A1(_02968_),
    .A2(_02978_),
    .B1(_02982_),
    .B2(_02799_),
    .X(_02986_));
 sky130_fd_sc_hd__o22ai_4 _08966_ (.A1(_02953_),
    .A2(_02954_),
    .B1(_02983_),
    .B2(_02985_),
    .Y(_02987_));
 sky130_fd_sc_hd__nor3_1 _08967_ (.A(_02953_),
    .B(_02954_),
    .C(_02985_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand3_2 _08968_ (.A(_02986_),
    .B(_02955_),
    .C(_02984_),
    .Y(_02989_));
 sky130_fd_sc_hd__o211ai_4 _08969_ (.A1(_02953_),
    .A2(_02954_),
    .B1(_02984_),
    .C1(_02986_),
    .Y(_02990_));
 sky130_fd_sc_hd__o21ai_2 _08970_ (.A1(_02983_),
    .A2(_02985_),
    .B1(_02955_),
    .Y(_02991_));
 sky130_fd_sc_hd__o2bb2ai_4 _08971_ (.A1_N(_02968_),
    .A2_N(_02971_),
    .B1(_02972_),
    .B2(_02974_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand4_4 _08972_ (.A(_02968_),
    .B(_02971_),
    .C(_02973_),
    .D(_02975_),
    .Y(_02994_));
 sky130_fd_sc_hd__o2bb2ai_1 _08973_ (.A1_N(_02968_),
    .A2_N(_02971_),
    .B1(_02976_),
    .B2(_02977_),
    .Y(_02995_));
 sky130_fd_sc_hd__a22oi_4 _08974_ (.A1(net30),
    .A2(net44),
    .B1(net33),
    .B2(net31),
    .Y(_02996_));
 sky130_fd_sc_hd__a22o_1 _08975_ (.A1(net30),
    .A2(net44),
    .B1(net33),
    .B2(net31),
    .X(_02997_));
 sky130_fd_sc_hd__and4_1 _08976_ (.A(net30),
    .B(net31),
    .C(net44),
    .D(net33),
    .X(_02998_));
 sky130_fd_sc_hd__nand4_2 _08977_ (.A(net30),
    .B(net31),
    .C(net44),
    .D(net33),
    .Y(_02999_));
 sky130_fd_sc_hd__nand2_1 _08978_ (.A(net29),
    .B(net55),
    .Y(_03000_));
 sky130_fd_sc_hd__o21ai_2 _08979_ (.A1(_03000_),
    .A2(_02996_),
    .B1(_02999_),
    .Y(_03001_));
 sky130_fd_sc_hd__o21a_2 _08980_ (.A1(_03000_),
    .A2(_02996_),
    .B1(_02999_),
    .X(_03002_));
 sky130_fd_sc_hd__o211ai_4 _08981_ (.A1(_00088_),
    .A2(_00341_),
    .B1(_02957_),
    .C1(_02960_),
    .Y(_03004_));
 sky130_fd_sc_hd__o21bai_4 _08982_ (.A1(_02956_),
    .A2(_02958_),
    .B1_N(_02961_),
    .Y(_03005_));
 sky130_fd_sc_hd__o22a_1 _08983_ (.A1(_00088_),
    .A2(_00341_),
    .B1(_02956_),
    .B2(_02958_),
    .X(_03006_));
 sky130_fd_sc_hd__a22o_1 _08984_ (.A1(net30),
    .A2(net55),
    .B1(_02957_),
    .B2(_02960_),
    .X(_03007_));
 sky130_fd_sc_hd__a41o_1 _08985_ (.A1(net32),
    .A2(net31),
    .A3(net44),
    .A4(net33),
    .B1(_02961_),
    .X(_03008_));
 sky130_fd_sc_hd__o21ai_2 _08986_ (.A1(_02956_),
    .A2(_03008_),
    .B1(_03001_),
    .Y(_03009_));
 sky130_fd_sc_hd__o211a_1 _08987_ (.A1(_02956_),
    .A2(_03008_),
    .B1(_03001_),
    .C1(_03007_),
    .X(_03010_));
 sky130_fd_sc_hd__o211ai_2 _08988_ (.A1(_02956_),
    .A2(_03008_),
    .B1(_03001_),
    .C1(_03007_),
    .Y(_03011_));
 sky130_fd_sc_hd__o211ai_4 _08989_ (.A1(_00077_),
    .A2(_00352_),
    .B1(_02898_),
    .C1(_02901_),
    .Y(_03012_));
 sky130_fd_sc_hd__o21bai_4 _08990_ (.A1(_02897_),
    .A2(_02900_),
    .B1_N(_02899_),
    .Y(_03013_));
 sky130_fd_sc_hd__o22a_1 _08991_ (.A1(_00077_),
    .A2(_00352_),
    .B1(_02897_),
    .B2(_02900_),
    .X(_03015_));
 sky130_fd_sc_hd__and4_1 _08992_ (.A(_02898_),
    .B(_02901_),
    .C(net27),
    .D(net60),
    .X(_03016_));
 sky130_fd_sc_hd__nand2_2 _08993_ (.A(_03012_),
    .B(_03013_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand3_4 _08994_ (.A(_03002_),
    .B(_03004_),
    .C(_03005_),
    .Y(_03018_));
 sky130_fd_sc_hd__a32oi_4 _08995_ (.A1(_03002_),
    .A2(_03004_),
    .A3(_03005_),
    .B1(_03012_),
    .B2(_03013_),
    .Y(_03019_));
 sky130_fd_sc_hd__a32o_1 _08996_ (.A1(_03002_),
    .A2(_03004_),
    .A3(_03005_),
    .B1(_03012_),
    .B2(_03013_),
    .X(_03020_));
 sky130_fd_sc_hd__a2bb2oi_4 _08997_ (.A1_N(_03006_),
    .A2_N(_03009_),
    .B1(_03017_),
    .B2(_03018_),
    .Y(_03021_));
 sky130_fd_sc_hd__a21oi_4 _08998_ (.A1(_02993_),
    .A2(_02994_),
    .B1(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__o221ai_2 _08999_ (.A1(_02969_),
    .A2(_02980_),
    .B1(_03010_),
    .B2(_03019_),
    .C1(_02995_),
    .Y(_03023_));
 sky130_fd_sc_hd__o21bai_4 _09000_ (.A1(_02913_),
    .A2(_02920_),
    .B1_N(_02919_),
    .Y(_03024_));
 sky130_fd_sc_hd__o21ai_1 _09001_ (.A1(_02913_),
    .A2(_02922_),
    .B1(_03024_),
    .Y(_03026_));
 sky130_fd_sc_hd__and3_1 _09002_ (.A(_02993_),
    .B(_03021_),
    .C(_02994_),
    .X(_03027_));
 sky130_fd_sc_hd__nand3_4 _09003_ (.A(_02993_),
    .B(_03021_),
    .C(_02994_),
    .Y(_03028_));
 sky130_fd_sc_hd__o211a_1 _09004_ (.A1(_02913_),
    .A2(_02922_),
    .B1(_03024_),
    .C1(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o211ai_2 _09005_ (.A1(_02913_),
    .A2(_02922_),
    .B1(_03024_),
    .C1(_03028_),
    .Y(_03030_));
 sky130_fd_sc_hd__a31oi_4 _09006_ (.A1(_02923_),
    .A2(_03024_),
    .A3(_03028_),
    .B1(_03022_),
    .Y(_03031_));
 sky130_fd_sc_hd__a31o_1 _09007_ (.A1(_02923_),
    .A2(_03024_),
    .A3(_03028_),
    .B1(_03022_),
    .X(_03032_));
 sky130_fd_sc_hd__o211a_1 _09008_ (.A1(_03022_),
    .A2(_03029_),
    .B1(_02987_),
    .C1(_02989_),
    .X(_03033_));
 sky130_fd_sc_hd__o211ai_4 _09009_ (.A1(_03022_),
    .A2(_03029_),
    .B1(_02987_),
    .C1(_02989_),
    .Y(_03034_));
 sky130_fd_sc_hd__and3b_1 _09010_ (.A_N(_02913_),
    .B(_02922_),
    .C(_02933_),
    .X(_03035_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_02933_),
    .B(_02924_),
    .Y(_03037_));
 sky130_fd_sc_hd__and3_1 _09012_ (.A(_02924_),
    .B(_02931_),
    .C(_02932_),
    .X(_03038_));
 sky130_fd_sc_hd__a21oi_1 _09013_ (.A1(_02931_),
    .A2(_02932_),
    .B1(_02924_),
    .Y(_03039_));
 sky130_fd_sc_hd__nor2_1 _09014_ (.A(_02934_),
    .B(_03035_),
    .Y(_03040_));
 sky130_fd_sc_hd__nor2_1 _09015_ (.A(_03038_),
    .B(_03039_),
    .Y(_03041_));
 sky130_fd_sc_hd__a21oi_1 _09016_ (.A1(_02987_),
    .A2(_02989_),
    .B1(_03032_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand3_2 _09017_ (.A(_02990_),
    .B(_02991_),
    .C(_03031_),
    .Y(_03043_));
 sky130_fd_sc_hd__a31oi_4 _09018_ (.A1(_03031_),
    .A2(_02991_),
    .A3(_02990_),
    .B1(_03041_),
    .Y(_03044_));
 sky130_fd_sc_hd__o211a_1 _09019_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_03043_),
    .C1(_03034_),
    .X(_03045_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_03044_),
    .B(_03034_),
    .Y(_03046_));
 sky130_fd_sc_hd__a21oi_1 _09021_ (.A1(_03043_),
    .A2(_03040_),
    .B1(_03033_),
    .Y(_03048_));
 sky130_fd_sc_hd__o2bb2a_1 _09022_ (.A1_N(_02936_),
    .A2_N(_02951_),
    .B1(_02949_),
    .B2(_02946_),
    .X(_03049_));
 sky130_fd_sc_hd__a2bb2o_1 _09023_ (.A1_N(_02946_),
    .A2_N(_02949_),
    .B1(_02951_),
    .B2(_02936_),
    .X(_03050_));
 sky130_fd_sc_hd__o21ai_1 _09024_ (.A1(_02835_),
    .A2(_02845_),
    .B1(_02848_),
    .Y(_03051_));
 sky130_fd_sc_hd__o221ai_2 _09025_ (.A1(_00033_),
    .A2(_00429_),
    .B1(_02835_),
    .B2(_02845_),
    .C1(_02848_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand3_1 _09026_ (.A(_03051_),
    .B(net36),
    .C(net1),
    .Y(_03053_));
 sky130_fd_sc_hd__o21ai_1 _09027_ (.A1(_00033_),
    .A2(_00429_),
    .B1(_03051_),
    .Y(_03054_));
 sky130_fd_sc_hd__o2111ai_2 _09028_ (.A1(_02835_),
    .A2(_02845_),
    .B1(_02848_),
    .C1(net36),
    .D1(net1),
    .Y(_03055_));
 sky130_fd_sc_hd__nand3_2 _09029_ (.A(_03053_),
    .B(_03049_),
    .C(_03052_),
    .Y(_03056_));
 sky130_fd_sc_hd__and3_1 _09030_ (.A(_03050_),
    .B(_03054_),
    .C(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__nand3_1 _09031_ (.A(_03050_),
    .B(_03054_),
    .C(_03055_),
    .Y(_03059_));
 sky130_fd_sc_hd__o2bb2a_1 _09032_ (.A1_N(_03056_),
    .A2_N(_03059_),
    .B1(_02927_),
    .B2(_02929_),
    .X(_03060_));
 sky130_fd_sc_hd__o2bb2ai_2 _09033_ (.A1_N(_03056_),
    .A2_N(_03059_),
    .B1(_02927_),
    .B2(_02929_),
    .Y(_03061_));
 sky130_fd_sc_hd__and3_1 _09034_ (.A(_03056_),
    .B(_03059_),
    .C(_02930_),
    .X(_03062_));
 sky130_fd_sc_hd__nand3_1 _09035_ (.A(_03056_),
    .B(_03059_),
    .C(_02930_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(_03061_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__o21bai_1 _09037_ (.A1(_02804_),
    .A2(_02808_),
    .B1_N(_02825_),
    .Y(_03065_));
 sky130_fd_sc_hd__o211ai_2 _09038_ (.A1(_02663_),
    .A2(_02807_),
    .B1(_02825_),
    .C1(_02806_),
    .Y(_03066_));
 sky130_fd_sc_hd__o221ai_4 _09039_ (.A1(_02663_),
    .A2(_02807_),
    .B1(_02823_),
    .B2(_02824_),
    .C1(_02806_),
    .Y(_03067_));
 sky130_fd_sc_hd__o21ai_2 _09040_ (.A1(_02804_),
    .A2(_02808_),
    .B1(_02825_),
    .Y(_03068_));
 sky130_fd_sc_hd__a21oi_1 _09041_ (.A1(_02986_),
    .A2(_02955_),
    .B1(_02983_),
    .Y(_03070_));
 sky130_fd_sc_hd__a21o_1 _09042_ (.A1(_02986_),
    .A2(_02955_),
    .B1(_02983_),
    .X(_03071_));
 sky130_fd_sc_hd__a2bb2oi_2 _09043_ (.A1_N(_02983_),
    .A2_N(_02988_),
    .B1(_03067_),
    .B2(_03068_),
    .Y(_03072_));
 sky130_fd_sc_hd__o211ai_2 _09044_ (.A1(_02983_),
    .A2(_02988_),
    .B1(_03065_),
    .C1(_03066_),
    .Y(_03073_));
 sky130_fd_sc_hd__a21oi_1 _09045_ (.A1(_03065_),
    .A2(_03066_),
    .B1(_03071_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand3_2 _09046_ (.A(_03067_),
    .B(_03068_),
    .C(_03070_),
    .Y(_03075_));
 sky130_fd_sc_hd__nor2_1 _09047_ (.A(_03064_),
    .B(_03074_),
    .Y(_03076_));
 sky130_fd_sc_hd__nand4_2 _09048_ (.A(_03061_),
    .B(_03063_),
    .C(_03073_),
    .D(_03075_),
    .Y(_03077_));
 sky130_fd_sc_hd__o22ai_2 _09049_ (.A1(_03060_),
    .A2(_03062_),
    .B1(_03072_),
    .B2(_03074_),
    .Y(_03078_));
 sky130_fd_sc_hd__o211ai_1 _09050_ (.A1(_03060_),
    .A2(_03062_),
    .B1(_03073_),
    .C1(_03075_),
    .Y(_03079_));
 sky130_fd_sc_hd__a21o_1 _09051_ (.A1(_03073_),
    .A2(_03075_),
    .B1(_03064_),
    .X(_03081_));
 sky130_fd_sc_hd__o211ai_4 _09052_ (.A1(_03033_),
    .A2(_03044_),
    .B1(_03077_),
    .C1(_03078_),
    .Y(_03082_));
 sky130_fd_sc_hd__nand3_1 _09053_ (.A(_03081_),
    .B(_03048_),
    .C(_03079_),
    .Y(_03083_));
 sky130_fd_sc_hd__a31oi_1 _09054_ (.A1(_03081_),
    .A2(_03048_),
    .A3(_03079_),
    .B1(_02935_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _09055_ (.A(_03084_),
    .B(_03082_),
    .Y(_03085_));
 sky130_fd_sc_hd__a2bb2oi_1 _09056_ (.A1_N(_02924_),
    .A2_N(_02933_),
    .B1(_03082_),
    .B2(_03083_),
    .Y(_03086_));
 sky130_fd_sc_hd__o2bb2ai_1 _09057_ (.A1_N(_03082_),
    .A2_N(_03083_),
    .B1(_02924_),
    .B2(_02933_),
    .Y(_03087_));
 sky130_fd_sc_hd__a21oi_1 _09058_ (.A1(_03082_),
    .A2(_03084_),
    .B1(_03086_),
    .Y(_03088_));
 sky130_fd_sc_hd__nand2_1 _09059_ (.A(_03085_),
    .B(_03087_),
    .Y(_03089_));
 sky130_fd_sc_hd__a22oi_4 _09060_ (.A1(net29),
    .A2(net44),
    .B1(net33),
    .B2(net30),
    .Y(_03090_));
 sky130_fd_sc_hd__a22o_1 _09061_ (.A1(net29),
    .A2(net44),
    .B1(net33),
    .B2(net30),
    .X(_03092_));
 sky130_fd_sc_hd__and4_1 _09062_ (.A(net30),
    .B(net29),
    .C(net44),
    .D(net33),
    .X(_03093_));
 sky130_fd_sc_hd__nand4_4 _09063_ (.A(net30),
    .B(net29),
    .C(net44),
    .D(net33),
    .Y(_03094_));
 sky130_fd_sc_hd__nand2_1 _09064_ (.A(net28),
    .B(net55),
    .Y(_03095_));
 sky130_fd_sc_hd__o21ai_4 _09065_ (.A1(_03095_),
    .A2(_03090_),
    .B1(_03094_),
    .Y(_03096_));
 sky130_fd_sc_hd__o211ai_1 _09066_ (.A1(_00099_),
    .A2(_00341_),
    .B1(_02997_),
    .C1(_02999_),
    .Y(_03097_));
 sky130_fd_sc_hd__o21bai_1 _09067_ (.A1(_02996_),
    .A2(_02998_),
    .B1_N(_03000_),
    .Y(_03098_));
 sky130_fd_sc_hd__o22a_1 _09068_ (.A1(_00099_),
    .A2(_00341_),
    .B1(_02996_),
    .B2(_02998_),
    .X(_03099_));
 sky130_fd_sc_hd__o21ai_2 _09069_ (.A1(_02996_),
    .A2(_02998_),
    .B1(_03000_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand4_2 _09070_ (.A(_02997_),
    .B(_02999_),
    .C(net29),
    .D(net55),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _09071_ (.A(_03096_),
    .B(_03101_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand3_4 _09072_ (.A(_03100_),
    .B(_03101_),
    .C(_03096_),
    .Y(_03104_));
 sky130_fd_sc_hd__a21oi_1 _09073_ (.A1(_03100_),
    .A2(_03101_),
    .B1(_03096_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand3b_2 _09074_ (.A_N(_03096_),
    .B(_03097_),
    .C(_03098_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(net26),
    .B(net60),
    .Y(_03107_));
 sky130_fd_sc_hd__and4_1 _09076_ (.A(net28),
    .B(net27),
    .C(net58),
    .D(net59),
    .X(_03108_));
 sky130_fd_sc_hd__nand4_1 _09077_ (.A(net28),
    .B(net27),
    .C(net58),
    .D(net59),
    .Y(_03109_));
 sky130_fd_sc_hd__a22oi_4 _09078_ (.A1(net28),
    .A2(net58),
    .B1(net59),
    .B2(net27),
    .Y(_03110_));
 sky130_fd_sc_hd__or2_1 _09079_ (.A(_03107_),
    .B(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__and4b_1 _09080_ (.A_N(_03110_),
    .B(net60),
    .C(net26),
    .D(_03109_),
    .X(_03112_));
 sky130_fd_sc_hd__o22a_1 _09081_ (.A1(_00044_),
    .A2(_00352_),
    .B1(_03108_),
    .B2(_03110_),
    .X(_03114_));
 sky130_fd_sc_hd__a2bb2o_1 _09082_ (.A1_N(_03108_),
    .A2_N(_03110_),
    .B1(net26),
    .B2(net60),
    .X(_03115_));
 sky130_fd_sc_hd__o21ai_1 _09083_ (.A1(_03108_),
    .A2(_03111_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__o2111ai_4 _09084_ (.A1(_03108_),
    .A2(_03111_),
    .B1(_03115_),
    .C1(_03106_),
    .D1(_03104_),
    .Y(_03117_));
 sky130_fd_sc_hd__o22a_1 _09085_ (.A1(_03099_),
    .A2(_03103_),
    .B1(_03105_),
    .B2(_03116_),
    .X(_03118_));
 sky130_fd_sc_hd__o211a_2 _09086_ (.A1(_03006_),
    .A2(_03009_),
    .B1(_03017_),
    .C1(_03018_),
    .X(_03119_));
 sky130_fd_sc_hd__a2bb2oi_4 _09087_ (.A1_N(_03015_),
    .A2_N(_03016_),
    .B1(_03018_),
    .B2(_03011_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21o_1 _09088_ (.A1(_03011_),
    .A2(_03018_),
    .B1(_03017_),
    .X(_03121_));
 sky130_fd_sc_hd__o21ai_1 _09089_ (.A1(_03010_),
    .A2(_03020_),
    .B1(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a21o_1 _09090_ (.A1(_03104_),
    .A2(_03117_),
    .B1(_03120_),
    .X(_03123_));
 sky130_fd_sc_hd__a211oi_4 _09091_ (.A1(_03104_),
    .A2(_03117_),
    .B1(_03119_),
    .C1(_03120_),
    .Y(_03125_));
 sky130_fd_sc_hd__a211o_1 _09092_ (.A1(_03104_),
    .A2(_03117_),
    .B1(_03119_),
    .C1(_03120_),
    .X(_03126_));
 sky130_fd_sc_hd__o221a_2 _09093_ (.A1(_03103_),
    .A2(_03099_),
    .B1(_03120_),
    .B2(_03119_),
    .C1(_03117_),
    .X(_03127_));
 sky130_fd_sc_hd__o21ai_1 _09094_ (.A1(_03119_),
    .A2(_03120_),
    .B1(_03118_),
    .Y(_03128_));
 sky130_fd_sc_hd__a22oi_4 _09095_ (.A1(net12),
    .A2(net62),
    .B1(net61),
    .B2(net23),
    .Y(_03129_));
 sky130_fd_sc_hd__a22o_1 _09096_ (.A1(net12),
    .A2(net62),
    .B1(net61),
    .B2(net23),
    .X(_03130_));
 sky130_fd_sc_hd__and4_1 _09097_ (.A(net12),
    .B(net23),
    .C(net62),
    .D(net61),
    .X(_03131_));
 sky130_fd_sc_hd__nand4_1 _09098_ (.A(net12),
    .B(net23),
    .C(net62),
    .D(net61),
    .Y(_03132_));
 sky130_fd_sc_hd__nand2_1 _09099_ (.A(net1),
    .B(net63),
    .Y(_03133_));
 sky130_fd_sc_hd__o41a_1 _09100_ (.A1(_00022_),
    .A2(_00055_),
    .A3(_00374_),
    .A4(_00385_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__a31o_1 _09101_ (.A1(_03130_),
    .A2(net63),
    .A3(net1),
    .B1(_03131_),
    .X(_03136_));
 sky130_fd_sc_hd__o2bb2ai_2 _09102_ (.A1_N(_02916_),
    .A2_N(_02917_),
    .B1(_00022_),
    .B2(_00396_),
    .Y(_03137_));
 sky130_fd_sc_hd__o21a_1 _09103_ (.A1(_00044_),
    .A2(_00352_),
    .B1(_03109_),
    .X(_03138_));
 sky130_fd_sc_hd__o21ai_1 _09104_ (.A1(_03107_),
    .A2(_03110_),
    .B1(_03109_),
    .Y(_03139_));
 sky130_fd_sc_hd__and3_1 _09105_ (.A(_02918_),
    .B(_03137_),
    .C(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__nand3_2 _09106_ (.A(_02918_),
    .B(_03137_),
    .C(_03139_),
    .Y(_03141_));
 sky130_fd_sc_hd__o2bb2a_1 _09107_ (.A1_N(_02918_),
    .A2_N(_03137_),
    .B1(_03138_),
    .B2(_03110_),
    .X(_03142_));
 sky130_fd_sc_hd__o2bb2ai_1 _09108_ (.A1_N(_02918_),
    .A2_N(_03137_),
    .B1(_03138_),
    .B2(_03110_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_2 _09109_ (.A(_03143_),
    .B(_03136_),
    .Y(_03144_));
 sky130_fd_sc_hd__a2bb2o_1 _09110_ (.A1_N(_03129_),
    .A2_N(_03134_),
    .B1(_03141_),
    .B2(_03143_),
    .X(_03145_));
 sky130_fd_sc_hd__o21a_1 _09111_ (.A1(_03140_),
    .A2(_03144_),
    .B1(_03145_),
    .X(_03147_));
 sky130_fd_sc_hd__o21ai_4 _09112_ (.A1(_03140_),
    .A2(_03144_),
    .B1(_03145_),
    .Y(_03148_));
 sky130_fd_sc_hd__a21oi_1 _09113_ (.A1(_03122_),
    .A2(_03118_),
    .B1(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__a21o_1 _09114_ (.A1(_03122_),
    .A2(_03118_),
    .B1(_03148_),
    .X(_03150_));
 sky130_fd_sc_hd__a21o_1 _09115_ (.A1(_03023_),
    .A2(_03028_),
    .B1(_03026_),
    .X(_03151_));
 sky130_fd_sc_hd__nand3_1 _09116_ (.A(_03023_),
    .B(_03026_),
    .C(_03028_),
    .Y(_03152_));
 sky130_fd_sc_hd__o21ai_1 _09117_ (.A1(_03022_),
    .A2(_03027_),
    .B1(_03026_),
    .Y(_03153_));
 sky130_fd_sc_hd__o221ai_4 _09118_ (.A1(_03022_),
    .A2(_03030_),
    .B1(_03125_),
    .B2(_03149_),
    .C1(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__a22o_1 _09119_ (.A1(net12),
    .A2(net64),
    .B1(net34),
    .B2(net1),
    .X(_03155_));
 sky130_fd_sc_hd__nand2_1 _09120_ (.A(_02927_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__o31a_1 _09121_ (.A1(_03129_),
    .A2(_03134_),
    .A3(_03142_),
    .B1(_03141_),
    .X(_03158_));
 sky130_fd_sc_hd__a21oi_2 _09122_ (.A1(_03141_),
    .A2(_03144_),
    .B1(_03156_),
    .Y(_03159_));
 sky130_fd_sc_hd__o311a_1 _09123_ (.A1(_03129_),
    .A2(_03134_),
    .A3(_03142_),
    .B1(_03156_),
    .C1(_03141_),
    .X(_03160_));
 sky130_fd_sc_hd__nor2_1 _09124_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__o2111ai_4 _09125_ (.A1(_03148_),
    .A2(_03127_),
    .B1(_03126_),
    .C1(_03152_),
    .D1(_03151_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand3_2 _09126_ (.A(_03154_),
    .B(_03161_),
    .C(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__a21boi_1 _09127_ (.A1(_03161_),
    .A2(_03162_),
    .B1_N(_03154_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_03154_),
    .B(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__a22oi_4 _09129_ (.A1(_02935_),
    .A2(_03037_),
    .B1(_03043_),
    .B2(_03034_),
    .Y(_03166_));
 sky130_fd_sc_hd__o22ai_1 _09130_ (.A1(_02934_),
    .A2(_03035_),
    .B1(_03042_),
    .B2(_03033_),
    .Y(_03167_));
 sky130_fd_sc_hd__a221oi_2 _09131_ (.A1(_03044_),
    .A2(_03034_),
    .B1(_03163_),
    .B2(_03154_),
    .C1(_03166_),
    .Y(_03169_));
 sky130_fd_sc_hd__a21oi_1 _09132_ (.A1(_03046_),
    .A2(_03167_),
    .B1(_03165_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21ai_1 _09133_ (.A1(_03045_),
    .A2(_03166_),
    .B1(_03164_),
    .Y(_03171_));
 sky130_fd_sc_hd__a21oi_1 _09134_ (.A1(_03171_),
    .A2(_03159_),
    .B1(_03169_),
    .Y(_03172_));
 sky130_fd_sc_hd__a32o_1 _09135_ (.A1(_03046_),
    .A2(_03165_),
    .A3(_03167_),
    .B1(_03171_),
    .B2(_03159_),
    .X(_03173_));
 sky130_fd_sc_hd__o311ai_2 _09136_ (.A1(_03045_),
    .A2(_03164_),
    .A3(_03166_),
    .B1(_03159_),
    .C1(_03171_),
    .Y(_03174_));
 sky130_fd_sc_hd__a21o_1 _09137_ (.A1(_03154_),
    .A2(_03162_),
    .B1(_03161_),
    .X(_03175_));
 sky130_fd_sc_hd__a22oi_2 _09138_ (.A1(net28),
    .A2(net44),
    .B1(net33),
    .B2(net29),
    .Y(_03176_));
 sky130_fd_sc_hd__a22o_1 _09139_ (.A1(net28),
    .A2(net44),
    .B1(net33),
    .B2(net29),
    .X(_03177_));
 sky130_fd_sc_hd__nand4_4 _09140_ (.A(net28),
    .B(net29),
    .C(net44),
    .D(net33),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _09141_ (.A(net27),
    .B(net55),
    .Y(_03180_));
 sky130_fd_sc_hd__o21ai_1 _09142_ (.A1(_03180_),
    .A2(_03176_),
    .B1(_03178_),
    .Y(_03181_));
 sky130_fd_sc_hd__o211ai_1 _09143_ (.A1(_00066_),
    .A2(_00341_),
    .B1(_03092_),
    .C1(_03094_),
    .Y(_03182_));
 sky130_fd_sc_hd__o21bai_1 _09144_ (.A1(_03090_),
    .A2(_03093_),
    .B1_N(_03095_),
    .Y(_03183_));
 sky130_fd_sc_hd__o22a_1 _09145_ (.A1(_00066_),
    .A2(_00341_),
    .B1(_03090_),
    .B2(_03093_),
    .X(_03184_));
 sky130_fd_sc_hd__a22o_1 _09146_ (.A1(net28),
    .A2(net55),
    .B1(_03092_),
    .B2(_03094_),
    .X(_03185_));
 sky130_fd_sc_hd__nand4_1 _09147_ (.A(_03092_),
    .B(_03094_),
    .C(net28),
    .D(net55),
    .Y(_03186_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_03181_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand3_1 _09149_ (.A(_03185_),
    .B(_03186_),
    .C(_03181_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand2_1 _09150_ (.A(net23),
    .B(net60),
    .Y(_03189_));
 sky130_fd_sc_hd__a22oi_1 _09151_ (.A1(net27),
    .A2(net58),
    .B1(net59),
    .B2(net26),
    .Y(_03191_));
 sky130_fd_sc_hd__a22o_1 _09152_ (.A1(net27),
    .A2(net58),
    .B1(net59),
    .B2(net26),
    .X(_03192_));
 sky130_fd_sc_hd__nand4_1 _09153_ (.A(net26),
    .B(net27),
    .C(net58),
    .D(net59),
    .Y(_03193_));
 sky130_fd_sc_hd__o211ai_1 _09154_ (.A1(_00055_),
    .A2(_00352_),
    .B1(_03192_),
    .C1(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__a21o_1 _09155_ (.A1(_03192_),
    .A2(_03193_),
    .B1(_03189_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_2 _09156_ (.A(_03194_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__nand3b_2 _09157_ (.A_N(_03181_),
    .B(_03182_),
    .C(_03183_),
    .Y(_03197_));
 sky130_fd_sc_hd__o211a_1 _09158_ (.A1(_03187_),
    .A2(_03184_),
    .B1(_03197_),
    .C1(_03196_),
    .X(_03198_));
 sky130_fd_sc_hd__o211ai_2 _09159_ (.A1(_03184_),
    .A2(_03187_),
    .B1(_03196_),
    .C1(_03197_),
    .Y(_03199_));
 sky130_fd_sc_hd__o2bb2ai_2 _09160_ (.A1_N(_03196_),
    .A2_N(_03197_),
    .B1(_03184_),
    .B2(_03187_),
    .Y(_03200_));
 sky130_fd_sc_hd__o2bb2ai_1 _09161_ (.A1_N(_03104_),
    .A2_N(_03106_),
    .B1(_03112_),
    .B2(_03114_),
    .Y(_03202_));
 sky130_fd_sc_hd__and3_1 _09162_ (.A(_03117_),
    .B(_03200_),
    .C(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__nand3_1 _09163_ (.A(_03117_),
    .B(_03200_),
    .C(_03202_),
    .Y(_03204_));
 sky130_fd_sc_hd__a21oi_1 _09164_ (.A1(_03117_),
    .A2(_03202_),
    .B1(_03200_),
    .Y(_03205_));
 sky130_fd_sc_hd__a21o_1 _09165_ (.A1(_03117_),
    .A2(_03202_),
    .B1(_03200_),
    .X(_03206_));
 sky130_fd_sc_hd__nand2_1 _09166_ (.A(net1),
    .B(net61),
    .Y(_03207_));
 sky130_fd_sc_hd__and4_2 _09167_ (.A(net12),
    .B(net1),
    .C(net62),
    .D(net61),
    .X(_03208_));
 sky130_fd_sc_hd__o21ai_1 _09168_ (.A1(_03189_),
    .A2(_03191_),
    .B1(_03193_),
    .Y(_03209_));
 sky130_fd_sc_hd__a211o_1 _09169_ (.A1(net1),
    .A2(net63),
    .B1(_03129_),
    .C1(_03131_),
    .X(_03210_));
 sky130_fd_sc_hd__a21o_1 _09170_ (.A1(_03130_),
    .A2(_03132_),
    .B1(_03133_),
    .X(_03211_));
 sky130_fd_sc_hd__a41o_1 _09171_ (.A1(net12),
    .A2(net23),
    .A3(net62),
    .A4(net61),
    .B1(_03133_),
    .X(_03213_));
 sky130_fd_sc_hd__a22o_1 _09172_ (.A1(net1),
    .A2(net63),
    .B1(_03130_),
    .B2(_03132_),
    .X(_03214_));
 sky130_fd_sc_hd__o211ai_1 _09173_ (.A1(_03129_),
    .A2(_03213_),
    .B1(_03209_),
    .C1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__nand3b_1 _09174_ (.A_N(_03209_),
    .B(_03210_),
    .C(_03211_),
    .Y(_03216_));
 sky130_fd_sc_hd__and3_1 _09175_ (.A(_03216_),
    .B(_03208_),
    .C(_03215_),
    .X(_03217_));
 sky130_fd_sc_hd__a21oi_1 _09176_ (.A1(_03215_),
    .A2(_03216_),
    .B1(_03208_),
    .Y(_03218_));
 sky130_fd_sc_hd__nor2_1 _09177_ (.A(_03217_),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__a21oi_1 _09178_ (.A1(_03219_),
    .A2(_03206_),
    .B1(_03203_),
    .Y(_03220_));
 sky130_fd_sc_hd__a21o_1 _09179_ (.A1(_03219_),
    .A2(_03206_),
    .B1(_03203_),
    .X(_03221_));
 sky130_fd_sc_hd__and3_1 _09180_ (.A(_03126_),
    .B(_03128_),
    .C(_03147_),
    .X(_03222_));
 sky130_fd_sc_hd__o21ai_1 _09181_ (.A1(_03125_),
    .A2(_03127_),
    .B1(_03148_),
    .Y(_03224_));
 sky130_fd_sc_hd__o211ai_1 _09182_ (.A1(_03119_),
    .A2(_03123_),
    .B1(_03128_),
    .C1(_03148_),
    .Y(_03225_));
 sky130_fd_sc_hd__o21ai_1 _09183_ (.A1(_03125_),
    .A2(_03127_),
    .B1(_03147_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(_03221_),
    .B(_03224_),
    .Y(_03227_));
 sky130_fd_sc_hd__o211ai_1 _09185_ (.A1(_03150_),
    .A2(_03125_),
    .B1(_03224_),
    .C1(_03221_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand3_1 _09186_ (.A(_03226_),
    .B(_03220_),
    .C(_03225_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21bo_1 _09187_ (.A1(_03216_),
    .A2(_03208_),
    .B1_N(_03215_),
    .X(_03230_));
 sky130_fd_sc_hd__and3_1 _09188_ (.A(_03230_),
    .B(net64),
    .C(net1),
    .X(_03231_));
 sky130_fd_sc_hd__a21o_1 _09189_ (.A1(net1),
    .A2(net64),
    .B1(_03230_),
    .X(_03232_));
 sky130_fd_sc_hd__and2b_1 _09190_ (.A_N(_03231_),
    .B(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__o2bb2ai_2 _09191_ (.A1_N(_03233_),
    .A2_N(_03229_),
    .B1(_03222_),
    .B2(_03227_),
    .Y(_03235_));
 sky130_fd_sc_hd__a21o_1 _09192_ (.A1(_03163_),
    .A2(_03175_),
    .B1(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__a31o_1 _09193_ (.A1(_03163_),
    .A2(_03175_),
    .A3(_03235_),
    .B1(_03231_),
    .X(_03237_));
 sky130_fd_sc_hd__o22ai_1 _09194_ (.A1(_03156_),
    .A2(_03158_),
    .B1(_03169_),
    .B2(_03170_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand4_1 _09195_ (.A(_03174_),
    .B(_03236_),
    .C(_03237_),
    .D(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__o21ai_1 _09196_ (.A1(_03172_),
    .A2(_03089_),
    .B1(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand4_1 _09197_ (.A(_03231_),
    .B(_03235_),
    .C(_03163_),
    .D(_03175_),
    .Y(_03241_));
 sky130_fd_sc_hd__o211ai_1 _09198_ (.A1(_03236_),
    .A2(_03231_),
    .B1(_03174_),
    .C1(_03238_),
    .Y(_03242_));
 sky130_fd_sc_hd__o2bb2ai_1 _09199_ (.A1_N(_03204_),
    .A2_N(_03206_),
    .B1(_03217_),
    .B2(_03218_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand3_1 _09200_ (.A(_03219_),
    .B(_03206_),
    .C(_03204_),
    .Y(_03244_));
 sky130_fd_sc_hd__o21ai_1 _09201_ (.A1(_03203_),
    .A2(_03205_),
    .B1(_03219_),
    .Y(_03246_));
 sky130_fd_sc_hd__o211ai_1 _09202_ (.A1(_03217_),
    .A2(_03218_),
    .B1(_03204_),
    .C1(_03206_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(net27),
    .B(net44),
    .Y(_03248_));
 sky130_fd_sc_hd__a22oi_4 _09204_ (.A1(net27),
    .A2(net44),
    .B1(net33),
    .B2(net28),
    .Y(_03249_));
 sky130_fd_sc_hd__and4_1 _09205_ (.A(net28),
    .B(net27),
    .C(net44),
    .D(net33),
    .X(_03250_));
 sky130_fd_sc_hd__nand4_2 _09206_ (.A(net28),
    .B(net27),
    .C(net44),
    .D(net33),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2_1 _09207_ (.A(net26),
    .B(net55),
    .Y(_03252_));
 sky130_fd_sc_hd__o21a_1 _09208_ (.A1(_00044_),
    .A2(_00341_),
    .B1(_03251_),
    .X(_03253_));
 sky130_fd_sc_hd__o21ai_1 _09209_ (.A1(_03252_),
    .A2(_03249_),
    .B1(_03251_),
    .Y(_03254_));
 sky130_fd_sc_hd__a22oi_4 _09210_ (.A1(net27),
    .A2(net55),
    .B1(_03177_),
    .B2(_03178_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand3_1 _09211_ (.A(_03178_),
    .B(net55),
    .C(net27),
    .Y(_03257_));
 sky130_fd_sc_hd__nor2_1 _09212_ (.A(_03176_),
    .B(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand4_1 _09213_ (.A(_03177_),
    .B(_03178_),
    .C(net27),
    .D(net55),
    .Y(_03259_));
 sky130_fd_sc_hd__o21ai_2 _09214_ (.A1(_03176_),
    .A2(_03257_),
    .B1(_03254_),
    .Y(_03260_));
 sky130_fd_sc_hd__nand3b_1 _09215_ (.A_N(_03255_),
    .B(_03259_),
    .C(_03254_),
    .Y(_03261_));
 sky130_fd_sc_hd__o22ai_4 _09216_ (.A1(_03249_),
    .A2(_03253_),
    .B1(_03255_),
    .B2(_03258_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(net12),
    .B(net60),
    .Y(_03263_));
 sky130_fd_sc_hd__and4_1 _09218_ (.A(net26),
    .B(net23),
    .C(net58),
    .D(net59),
    .X(_03264_));
 sky130_fd_sc_hd__nand4_1 _09219_ (.A(net26),
    .B(net23),
    .C(net58),
    .D(net59),
    .Y(_03265_));
 sky130_fd_sc_hd__a22o_1 _09220_ (.A1(net26),
    .A2(net58),
    .B1(net59),
    .B2(net23),
    .X(_03266_));
 sky130_fd_sc_hd__and4_1 _09221_ (.A(_03266_),
    .B(net60),
    .C(net12),
    .D(_03265_),
    .X(_03268_));
 sky130_fd_sc_hd__o2bb2a_1 _09222_ (.A1_N(_03265_),
    .A2_N(_03266_),
    .B1(_00022_),
    .B2(_00352_),
    .X(_03269_));
 sky130_fd_sc_hd__a21o_1 _09223_ (.A1(_03265_),
    .A2(_03266_),
    .B1(_03263_),
    .X(_03270_));
 sky130_fd_sc_hd__o211ai_1 _09224_ (.A1(_00022_),
    .A2(_00352_),
    .B1(_03265_),
    .C1(_03266_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _09225_ (.A(_03270_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__o2bb2ai_2 _09226_ (.A1_N(_03272_),
    .A2_N(_03262_),
    .B1(_03260_),
    .B2(_03255_),
    .Y(_03273_));
 sky130_fd_sc_hd__a21oi_1 _09227_ (.A1(_03188_),
    .A2(_03197_),
    .B1(_03196_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21o_1 _09228_ (.A1(_03188_),
    .A2(_03197_),
    .B1(_03196_),
    .X(_03275_));
 sky130_fd_sc_hd__o21bai_2 _09229_ (.A1(_03198_),
    .A2(_03274_),
    .B1_N(_03273_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand3_2 _09230_ (.A(_03199_),
    .B(_03273_),
    .C(_03275_),
    .Y(_03277_));
 sky130_fd_sc_hd__o22a_1 _09231_ (.A1(_00033_),
    .A2(_00374_),
    .B1(_00385_),
    .B2(_00022_),
    .X(_03279_));
 sky130_fd_sc_hd__or2_1 _09232_ (.A(_03208_),
    .B(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__a31o_1 _09233_ (.A1(_03266_),
    .A2(net60),
    .A3(net12),
    .B1(_03264_),
    .X(_03281_));
 sky130_fd_sc_hd__inv_2 _09234_ (.A(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__nor3b_2 _09235_ (.A(_03208_),
    .B(_03279_),
    .C_N(_03281_),
    .Y(_03283_));
 sky130_fd_sc_hd__o21a_1 _09236_ (.A1(_03208_),
    .A2(_03279_),
    .B1(_03282_),
    .X(_03284_));
 sky130_fd_sc_hd__nor2_1 _09237_ (.A(_03283_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__a31o_1 _09238_ (.A1(_03199_),
    .A2(_03273_),
    .A3(_03275_),
    .B1(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__a21boi_1 _09239_ (.A1(_03276_),
    .A2(_03285_),
    .B1_N(_03277_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand4_1 _09240_ (.A(_03243_),
    .B(_03244_),
    .C(_03276_),
    .D(_03286_),
    .Y(_03288_));
 sky130_fd_sc_hd__nand3_1 _09241_ (.A(_03246_),
    .B(_03247_),
    .C(_03287_),
    .Y(_03290_));
 sky130_fd_sc_hd__a21boi_1 _09242_ (.A1(_03290_),
    .A2(_03283_),
    .B1_N(_03288_),
    .Y(_03291_));
 sky130_fd_sc_hd__and3_1 _09243_ (.A(_03228_),
    .B(_03229_),
    .C(_03233_),
    .X(_03292_));
 sky130_fd_sc_hd__a21oi_1 _09244_ (.A1(_03228_),
    .A2(_03229_),
    .B1(_03233_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor3_1 _09245_ (.A(_03291_),
    .B(_03292_),
    .C(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__o21ai_1 _09246_ (.A1(_03292_),
    .A2(_03293_),
    .B1(_03291_),
    .Y(_03295_));
 sky130_fd_sc_hd__o2bb2ai_1 _09247_ (.A1_N(_03288_),
    .A2_N(_03290_),
    .B1(_03280_),
    .B2(_03282_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand3_1 _09248_ (.A(_03290_),
    .B(_03283_),
    .C(_03288_),
    .Y(_03297_));
 sky130_fd_sc_hd__a22o_2 _09249_ (.A1(net26),
    .A2(net44),
    .B1(net33),
    .B2(net27),
    .X(_03298_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(net26),
    .B(net33),
    .Y(_03299_));
 sky130_fd_sc_hd__nand4_2 _09251_ (.A(net26),
    .B(net27),
    .C(net44),
    .D(net33),
    .Y(_03301_));
 sky130_fd_sc_hd__o21ai_2 _09252_ (.A1(_00055_),
    .A2(_00341_),
    .B1(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand3_1 _09253_ (.A(_03251_),
    .B(net55),
    .C(net26),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _09254_ (.A(_03249_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand4b_1 _09255_ (.A_N(_03249_),
    .B(_03251_),
    .C(net26),
    .D(net55),
    .Y(_03305_));
 sky130_fd_sc_hd__o22a_1 _09256_ (.A1(_00044_),
    .A2(_00341_),
    .B1(_03249_),
    .B2(_03250_),
    .X(_03306_));
 sky130_fd_sc_hd__o21ai_1 _09257_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_03252_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand4_2 _09258_ (.A(_03298_),
    .B(_03302_),
    .C(_03305_),
    .D(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__a22oi_1 _09259_ (.A1(_03298_),
    .A2(_03302_),
    .B1(_03305_),
    .B2(_03307_),
    .Y(_03309_));
 sky130_fd_sc_hd__o2bb2ai_1 _09260_ (.A1_N(_03298_),
    .A2_N(_03302_),
    .B1(_03304_),
    .B2(_03306_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(net12),
    .B(net59),
    .Y(_03312_));
 sky130_fd_sc_hd__a22o_1 _09262_ (.A1(net23),
    .A2(net58),
    .B1(net59),
    .B2(net12),
    .X(_03313_));
 sky130_fd_sc_hd__nand4_2 _09263_ (.A(net12),
    .B(net23),
    .C(net58),
    .D(net59),
    .Y(_03314_));
 sky130_fd_sc_hd__o2bb2a_1 _09264_ (.A1_N(_03313_),
    .A2_N(_03314_),
    .B1(_00033_),
    .B2(_00352_),
    .X(_03315_));
 sky130_fd_sc_hd__a22o_1 _09265_ (.A1(net1),
    .A2(net60),
    .B1(_03313_),
    .B2(_03314_),
    .X(_03316_));
 sky130_fd_sc_hd__and4_1 _09266_ (.A(_03313_),
    .B(_03314_),
    .C(net1),
    .D(net60),
    .X(_03317_));
 sky130_fd_sc_hd__nand4_2 _09267_ (.A(_03313_),
    .B(_03314_),
    .C(net1),
    .D(net60),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(_03316_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__o21a_1 _09269_ (.A1(_03319_),
    .A2(_03309_),
    .B1(_03308_),
    .X(_03320_));
 sky130_fd_sc_hd__o21ai_1 _09270_ (.A1(_03319_),
    .A2(_03309_),
    .B1(_03308_),
    .Y(_03321_));
 sky130_fd_sc_hd__o211ai_1 _09271_ (.A1(_03255_),
    .A2(_03260_),
    .B1(_03262_),
    .C1(_03272_),
    .Y(_03323_));
 sky130_fd_sc_hd__o2bb2ai_1 _09272_ (.A1_N(_03261_),
    .A2_N(_03262_),
    .B1(_03268_),
    .B2(_03269_),
    .Y(_03324_));
 sky130_fd_sc_hd__o221ai_2 _09273_ (.A1(_03255_),
    .A2(_03260_),
    .B1(_03268_),
    .B2(_03269_),
    .C1(_03262_),
    .Y(_03325_));
 sky130_fd_sc_hd__a22o_1 _09274_ (.A1(_03261_),
    .A2(_03262_),
    .B1(_03270_),
    .B2(_03271_),
    .X(_03326_));
 sky130_fd_sc_hd__nand3_1 _09275_ (.A(_03321_),
    .B(_03323_),
    .C(_03324_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand3_2 _09276_ (.A(_03326_),
    .B(_03320_),
    .C(_03325_),
    .Y(_03328_));
 sky130_fd_sc_hd__o31a_1 _09277_ (.A1(_00055_),
    .A2(_00330_),
    .A3(_03312_),
    .B1(_03318_),
    .X(_03329_));
 sky130_fd_sc_hd__a21oi_1 _09278_ (.A1(_03314_),
    .A2(_03318_),
    .B1(_03207_),
    .Y(_03330_));
 sky130_fd_sc_hd__or3_1 _09279_ (.A(_00033_),
    .B(_00385_),
    .C(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__o311a_1 _09280_ (.A1(_00055_),
    .A2(_00330_),
    .A3(_03312_),
    .B1(_03318_),
    .C1(_03207_),
    .X(_03332_));
 sky130_fd_sc_hd__nor2_1 _09281_ (.A(_03330_),
    .B(_03332_),
    .Y(_03334_));
 sky130_fd_sc_hd__a21boi_1 _09282_ (.A1(_03328_),
    .A2(_03334_),
    .B1_N(_03327_),
    .Y(_03335_));
 sky130_fd_sc_hd__a21bo_1 _09283_ (.A1(_03328_),
    .A2(_03334_),
    .B1_N(_03327_),
    .X(_03336_));
 sky130_fd_sc_hd__a21bo_1 _09284_ (.A1(_03276_),
    .A2(_03277_),
    .B1_N(_03285_),
    .X(_03337_));
 sky130_fd_sc_hd__o211ai_1 _09285_ (.A1(_03283_),
    .A2(_03284_),
    .B1(_03276_),
    .C1(_03277_),
    .Y(_03338_));
 sky130_fd_sc_hd__o2bb2ai_1 _09286_ (.A1_N(_03276_),
    .A2_N(_03277_),
    .B1(_03283_),
    .B2(_03284_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand3_1 _09287_ (.A(_03276_),
    .B(_03277_),
    .C(_03285_),
    .Y(_03340_));
 sky130_fd_sc_hd__and3_1 _09288_ (.A(_03336_),
    .B(_03339_),
    .C(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__nand3_1 _09289_ (.A(_03336_),
    .B(_03339_),
    .C(_03340_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand3_1 _09290_ (.A(_03337_),
    .B(_03338_),
    .C(_03335_),
    .Y(_03343_));
 sky130_fd_sc_hd__a31oi_1 _09291_ (.A1(_03337_),
    .A2(_03338_),
    .A3(_03335_),
    .B1(_03331_),
    .Y(_03345_));
 sky130_fd_sc_hd__o211ai_1 _09292_ (.A1(_03341_),
    .A2(_03345_),
    .B1(_03296_),
    .C1(_03297_),
    .Y(_03346_));
 sky130_fd_sc_hd__a211o_1 _09293_ (.A1(_03296_),
    .A2(_03297_),
    .B1(_03341_),
    .C1(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__o2bb2ai_1 _09294_ (.A1_N(_03342_),
    .A2_N(_03343_),
    .B1(_03207_),
    .B2(_03329_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand4_4 _09295_ (.A(net26),
    .B(net23),
    .C(net44),
    .D(net33),
    .Y(_03349_));
 sky130_fd_sc_hd__a22o_1 _09296_ (.A1(net23),
    .A2(net44),
    .B1(net33),
    .B2(net26),
    .X(_03350_));
 sky130_fd_sc_hd__nand4_4 _09297_ (.A(_03350_),
    .B(net55),
    .C(net12),
    .D(_03349_),
    .Y(_03351_));
 sky130_fd_sc_hd__a22oi_2 _09298_ (.A1(net23),
    .A2(net55),
    .B1(_03298_),
    .B2(_03301_),
    .Y(_03352_));
 sky130_fd_sc_hd__o2111a_1 _09299_ (.A1(_03248_),
    .A2(_03299_),
    .B1(net23),
    .C1(net55),
    .D1(_03298_),
    .X(_03353_));
 sky130_fd_sc_hd__a21o_1 _09300_ (.A1(_03349_),
    .A2(_03351_),
    .B1(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__a211o_1 _09301_ (.A1(_03349_),
    .A2(_03351_),
    .B1(_03352_),
    .C1(_03353_),
    .X(_03356_));
 sky130_fd_sc_hd__o211ai_2 _09302_ (.A1(_03352_),
    .A2(_03353_),
    .B1(_03349_),
    .C1(_03351_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_1 _09303_ (.A(net1),
    .B(net58),
    .Y(_03358_));
 sky130_fd_sc_hd__or4_1 _09304_ (.A(_00022_),
    .B(_00033_),
    .C(_00330_),
    .D(_00363_),
    .X(_03359_));
 sky130_fd_sc_hd__a22o_1 _09305_ (.A1(net12),
    .A2(net58),
    .B1(net59),
    .B2(net1),
    .X(_03360_));
 sky130_fd_sc_hd__o31a_1 _09306_ (.A1(_00022_),
    .A2(_00363_),
    .A3(_03358_),
    .B1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__o2111ai_1 _09307_ (.A1(_03312_),
    .A2(_03358_),
    .B1(_03360_),
    .C1(_03356_),
    .D1(_03357_),
    .Y(_03362_));
 sky130_fd_sc_hd__o2bb2ai_1 _09308_ (.A1_N(_03361_),
    .A2_N(_03357_),
    .B1(_03354_),
    .B2(_03352_),
    .Y(_03363_));
 sky130_fd_sc_hd__o2bb2ai_1 _09309_ (.A1_N(_03308_),
    .A2_N(_03310_),
    .B1(_03315_),
    .B2(_03317_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand4_1 _09310_ (.A(_03308_),
    .B(_03310_),
    .C(_03316_),
    .D(_03318_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand3_1 _09311_ (.A(_03363_),
    .B(_03364_),
    .C(_03365_),
    .Y(_03367_));
 sky130_fd_sc_hd__and3_1 _09312_ (.A(_03327_),
    .B(_03328_),
    .C(_03334_),
    .X(_03368_));
 sky130_fd_sc_hd__nand3_1 _09313_ (.A(_03327_),
    .B(_03328_),
    .C(_03334_),
    .Y(_03369_));
 sky130_fd_sc_hd__o2bb2ai_1 _09314_ (.A1_N(_03327_),
    .A2_N(_03328_),
    .B1(_03330_),
    .B2(_03332_),
    .Y(_03370_));
 sky130_fd_sc_hd__a21oi_1 _09315_ (.A1(_03364_),
    .A2(_03365_),
    .B1(_03363_),
    .Y(_03371_));
 sky130_fd_sc_hd__a21o_1 _09316_ (.A1(_03364_),
    .A2(_03365_),
    .B1(_03363_),
    .X(_03372_));
 sky130_fd_sc_hd__o2bb2ai_1 _09317_ (.A1_N(_03367_),
    .A2_N(_03372_),
    .B1(_03312_),
    .B2(_03358_),
    .Y(_03373_));
 sky130_fd_sc_hd__a22o_1 _09318_ (.A1(_03356_),
    .A2(_03357_),
    .B1(_03359_),
    .B2(_03360_),
    .X(_03374_));
 sky130_fd_sc_hd__a22o_1 _09319_ (.A1(net12),
    .A2(net55),
    .B1(_03349_),
    .B2(_03350_),
    .X(_03375_));
 sky130_fd_sc_hd__and2_1 _09320_ (.A(net1),
    .B(net55),
    .X(_03376_));
 sky130_fd_sc_hd__a22o_1 _09321_ (.A1(net12),
    .A2(net44),
    .B1(net33),
    .B2(net23),
    .X(_03378_));
 sky130_fd_sc_hd__and4_1 _09322_ (.A(net12),
    .B(net23),
    .C(net44),
    .D(net33),
    .X(_03379_));
 sky130_fd_sc_hd__a31o_1 _09323_ (.A1(_03378_),
    .A2(net55),
    .A3(net1),
    .B1(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__nand4_1 _09324_ (.A(net12),
    .B(net1),
    .C(net44),
    .D(net33),
    .Y(_03381_));
 sky130_fd_sc_hd__a21oi_1 _09325_ (.A1(_00055_),
    .A2(net55),
    .B1(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__o31a_1 _09326_ (.A1(_00055_),
    .A2(_00319_),
    .A3(_03376_),
    .B1(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__and4_1 _09327_ (.A(net1),
    .B(net58),
    .C(_03380_),
    .D(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__a32o_1 _09328_ (.A1(_03351_),
    .A2(_03384_),
    .A3(_03375_),
    .B1(_03374_),
    .B2(_03362_),
    .X(_03385_));
 sky130_fd_sc_hd__a21o_1 _09329_ (.A1(net1),
    .A2(net58),
    .B1(_03383_),
    .X(_03386_));
 sky130_fd_sc_hd__a32o_1 _09330_ (.A1(net1),
    .A2(net58),
    .A3(_03383_),
    .B1(_03375_),
    .B2(_03351_),
    .X(_03387_));
 sky130_fd_sc_hd__o21a_1 _09331_ (.A1(_03380_),
    .A2(_03386_),
    .B1(_03387_),
    .X(_03389_));
 sky130_fd_sc_hd__a21o_1 _09332_ (.A1(_03380_),
    .A2(_03386_),
    .B1(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__o21ai_1 _09333_ (.A1(_03359_),
    .A2(_03371_),
    .B1(_03367_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _09334_ (.A(_03370_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21oi_1 _09335_ (.A1(_03369_),
    .A2(_03370_),
    .B1(_03391_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand3b_1 _09336_ (.A_N(_03359_),
    .B(_03367_),
    .C(_03372_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand4_1 _09337_ (.A(_03373_),
    .B(_03385_),
    .C(_03390_),
    .D(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__o22ai_1 _09338_ (.A1(_03368_),
    .A2(_03392_),
    .B1(_03395_),
    .B2(_03393_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand3_1 _09339_ (.A(_03342_),
    .B(_03343_),
    .C(_03330_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand3_1 _09340_ (.A(_03348_),
    .B(_03396_),
    .C(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03346_),
    .B(_03398_),
    .Y(_03400_));
 sky130_fd_sc_hd__a31oi_2 _09342_ (.A1(_03295_),
    .A2(_03347_),
    .A3(_03400_),
    .B1(_03294_),
    .Y(_03401_));
 sky130_fd_sc_hd__a21oi_1 _09343_ (.A1(_03241_),
    .A2(_03242_),
    .B1(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__a21boi_1 _09344_ (.A1(_03083_),
    .A2(_02934_),
    .B1_N(_03082_),
    .Y(_03403_));
 sky130_fd_sc_hd__a21oi_1 _09345_ (.A1(_02930_),
    .A2(_03056_),
    .B1(_03057_),
    .Y(_03404_));
 sky130_fd_sc_hd__o22ai_2 _09346_ (.A1(_02859_),
    .A2(_02862_),
    .B1(_02865_),
    .B2(_02833_),
    .Y(_03405_));
 sky130_fd_sc_hd__a31o_1 _09347_ (.A1(_03061_),
    .A2(_03063_),
    .A3(_03075_),
    .B1(_03072_),
    .X(_03406_));
 sky130_fd_sc_hd__o211a_1 _09348_ (.A1(_03072_),
    .A2(_03076_),
    .B1(_03405_),
    .C1(_02867_),
    .X(_03407_));
 sky130_fd_sc_hd__o211ai_1 _09349_ (.A1(_03072_),
    .A2(_03076_),
    .B1(_03405_),
    .C1(_02867_),
    .Y(_03408_));
 sky130_fd_sc_hd__a21oi_1 _09350_ (.A1(_02867_),
    .A2(_03405_),
    .B1(_03406_),
    .Y(_03409_));
 sky130_fd_sc_hd__a21o_1 _09351_ (.A1(_02867_),
    .A2(_03405_),
    .B1(_03406_),
    .X(_03411_));
 sky130_fd_sc_hd__nand3_1 _09352_ (.A(_03411_),
    .B(_03404_),
    .C(_03408_),
    .Y(_03412_));
 sky130_fd_sc_hd__o22ai_1 _09353_ (.A1(_03057_),
    .A2(_03062_),
    .B1(_03407_),
    .B2(_03409_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand3_1 _09354_ (.A(_03413_),
    .B(_03403_),
    .C(_03412_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_1 _09355_ (.A1(_03173_),
    .A2(_03088_),
    .B1(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__o21bai_2 _09356_ (.A1(_03240_),
    .A2(_03402_),
    .B1_N(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21a_1 _09357_ (.A1(_03404_),
    .A2(_03409_),
    .B1(_03408_),
    .X(_03417_));
 sky130_fd_sc_hd__nand3_1 _09358_ (.A(_02875_),
    .B(_02876_),
    .C(_02879_),
    .Y(_03418_));
 sky130_fd_sc_hd__a21o_1 _09359_ (.A1(_02875_),
    .A2(_02876_),
    .B1(_02879_),
    .X(_03419_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__a22o_1 _09361_ (.A1(_03082_),
    .A2(_03085_),
    .B1(_03412_),
    .B2(_03413_),
    .X(_03422_));
 sky130_fd_sc_hd__o211ai_4 _09362_ (.A1(_03417_),
    .A2(_03420_),
    .B1(_03422_),
    .C1(_03416_),
    .Y(_03423_));
 sky130_fd_sc_hd__o2bb2ai_1 _09363_ (.A1_N(_02888_),
    .A2_N(_02895_),
    .B1(_02715_),
    .B2(_02878_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand2_1 _09364_ (.A(_03417_),
    .B(_03420_),
    .Y(_03425_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_03424_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_02769_),
    .B(_02896_),
    .Y(_03427_));
 sky130_fd_sc_hd__a31oi_1 _09367_ (.A1(_02888_),
    .A2(_02891_),
    .A3(_02892_),
    .B1(_03426_),
    .Y(_03428_));
 sky130_fd_sc_hd__a21oi_2 _09368_ (.A1(_03428_),
    .A2(_03423_),
    .B1(_03427_),
    .Y(_03429_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(_02637_),
    .B(_02566_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21o_1 _09370_ (.A1(_02565_),
    .A2(_02638_),
    .B1(_02768_),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_1 _09371_ (.A(_03430_),
    .B(_03431_),
    .Y(_03433_));
 sky130_fd_sc_hd__o22ai_4 _09372_ (.A1(_02566_),
    .A2(_02637_),
    .B1(_03433_),
    .B2(_03429_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21boi_1 _09373_ (.A1(_02633_),
    .A2(_02634_),
    .B1_N(_02632_),
    .Y(_03435_));
 sky130_fd_sc_hd__a2bb2o_1 _09374_ (.A1_N(_02580_),
    .A2_N(_02586_),
    .B1(_02584_),
    .B2(_02568_),
    .X(_03436_));
 sky130_fd_sc_hd__a21oi_1 _09375_ (.A1(_02592_),
    .A2(_02626_),
    .B1(_02623_),
    .Y(_03437_));
 sky130_fd_sc_hd__a21o_1 _09376_ (.A1(_02592_),
    .A2(_02626_),
    .B1(_02623_),
    .X(_03438_));
 sky130_fd_sc_hd__o22a_1 _09377_ (.A1(_02595_),
    .A2(_02603_),
    .B1(_02606_),
    .B2(_02601_),
    .X(_03439_));
 sky130_fd_sc_hd__o21ai_1 _09378_ (.A1(_02601_),
    .A2(_02606_),
    .B1(_02605_),
    .Y(_03440_));
 sky130_fd_sc_hd__o2bb2ai_1 _09379_ (.A1_N(_02055_),
    .A2_N(_02056_),
    .B1(_02059_),
    .B2(_02060_),
    .Y(_03441_));
 sky130_fd_sc_hd__o211ai_1 _09380_ (.A1(_01852_),
    .A2(_02058_),
    .B1(_02056_),
    .C1(_02055_),
    .Y(_03442_));
 sky130_fd_sc_hd__o2bb2ai_1 _09381_ (.A1_N(_02055_),
    .A2_N(_02056_),
    .B1(_02058_),
    .B2(_01852_),
    .Y(_03444_));
 sky130_fd_sc_hd__o211ai_1 _09382_ (.A1(_02059_),
    .A2(_02060_),
    .B1(_02055_),
    .C1(_02056_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand3_2 _09383_ (.A(_03439_),
    .B(_03441_),
    .C(_03442_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand3_2 _09384_ (.A(_03440_),
    .B(_03444_),
    .C(_03445_),
    .Y(_03447_));
 sky130_fd_sc_hd__o32a_1 _09385_ (.A1(_02049_),
    .A2(_02569_),
    .A3(_02572_),
    .B1(_00473_),
    .B2(_00033_),
    .X(_03448_));
 sky130_fd_sc_hd__o21ai_1 _09386_ (.A1(_01851_),
    .A2(_02575_),
    .B1(_02576_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand3_2 _09387_ (.A(_03446_),
    .B(_03447_),
    .C(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__o2bb2ai_2 _09388_ (.A1_N(_03446_),
    .A2_N(_03447_),
    .B1(_03448_),
    .B2(_02575_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(_03450_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__o21ai_2 _09390_ (.A1(_02614_),
    .A2(_02610_),
    .B1(_02617_),
    .Y(_03453_));
 sky130_fd_sc_hd__o21a_1 _09391_ (.A1(_02614_),
    .A2(_02610_),
    .B1(_02617_),
    .X(_03455_));
 sky130_fd_sc_hd__o211ai_2 _09392_ (.A1(_02007_),
    .A2(_02008_),
    .B1(_01974_),
    .C1(_01977_),
    .Y(_03456_));
 sky130_fd_sc_hd__o2bb2ai_1 _09393_ (.A1_N(_01974_),
    .A2_N(_01977_),
    .B1(_02009_),
    .B2(_02011_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand3_2 _09394_ (.A(_01974_),
    .B(_01977_),
    .C(_02014_),
    .Y(_03458_));
 sky130_fd_sc_hd__o2bb2ai_2 _09395_ (.A1_N(_01974_),
    .A2_N(_01977_),
    .B1(_02007_),
    .B2(_02008_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand3_2 _09396_ (.A(_03457_),
    .B(_03453_),
    .C(_03456_),
    .Y(_03460_));
 sky130_fd_sc_hd__and3_1 _09397_ (.A(_03455_),
    .B(_03458_),
    .C(_03459_),
    .X(_03461_));
 sky130_fd_sc_hd__o2111ai_4 _09398_ (.A1(_02610_),
    .A2(_02614_),
    .B1(_02617_),
    .C1(_03458_),
    .D1(_03459_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand3_1 _09399_ (.A(_03452_),
    .B(_03460_),
    .C(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__a21o_1 _09400_ (.A1(_03460_),
    .A2(_03462_),
    .B1(_03452_),
    .X(_03464_));
 sky130_fd_sc_hd__nand4_1 _09401_ (.A(_03450_),
    .B(_03451_),
    .C(_03460_),
    .D(_03462_),
    .Y(_03466_));
 sky130_fd_sc_hd__a22o_1 _09402_ (.A1(_03450_),
    .A2(_03451_),
    .B1(_03460_),
    .B2(_03462_),
    .X(_03467_));
 sky130_fd_sc_hd__nand3_1 _09403_ (.A(_03438_),
    .B(_03466_),
    .C(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand3_1 _09404_ (.A(_03464_),
    .B(_03437_),
    .C(_03463_),
    .Y(_03469_));
 sky130_fd_sc_hd__nand3_1 _09405_ (.A(_03468_),
    .B(_03469_),
    .C(_03436_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21o_1 _09406_ (.A1(_03468_),
    .A2(_03469_),
    .B1(_03436_),
    .X(_03471_));
 sky130_fd_sc_hd__nand3_1 _09407_ (.A(_03435_),
    .B(_03470_),
    .C(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__a32o_1 _09408_ (.A1(_03438_),
    .A2(_03466_),
    .A3(_03467_),
    .B1(_03469_),
    .B2(_03436_),
    .X(_03473_));
 sky130_fd_sc_hd__a21bo_1 _09409_ (.A1(_03446_),
    .A2(_03449_),
    .B1_N(_03447_),
    .X(_03474_));
 sky130_fd_sc_hd__a32oi_2 _09410_ (.A1(_03457_),
    .A2(_03453_),
    .A3(_03456_),
    .B1(_03451_),
    .B2(_03450_),
    .Y(_03475_));
 sky130_fd_sc_hd__a32oi_1 _09411_ (.A1(_03455_),
    .A2(_03458_),
    .A3(_03459_),
    .B1(_03460_),
    .B2(_03452_),
    .Y(_03477_));
 sky130_fd_sc_hd__nand3_1 _09412_ (.A(_02022_),
    .B(_02025_),
    .C(_02075_),
    .Y(_03478_));
 sky130_fd_sc_hd__o21bai_1 _09413_ (.A1(_02021_),
    .A2(_02023_),
    .B1_N(_02075_),
    .Y(_03479_));
 sky130_fd_sc_hd__o2111ai_1 _09414_ (.A1(_02070_),
    .A2(_02073_),
    .B1(_02074_),
    .C1(_02025_),
    .D1(_02022_),
    .Y(_03480_));
 sky130_fd_sc_hd__o21ai_1 _09415_ (.A1(_02021_),
    .A2(_02023_),
    .B1(_02075_),
    .Y(_03481_));
 sky130_fd_sc_hd__o211ai_2 _09416_ (.A1(_03461_),
    .A2(_03475_),
    .B1(_03478_),
    .C1(_03479_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand3_1 _09417_ (.A(_03481_),
    .B(_03477_),
    .C(_03480_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand3_1 _09418_ (.A(_03482_),
    .B(_03483_),
    .C(_03474_),
    .Y(_03484_));
 sky130_fd_sc_hd__a21o_1 _09419_ (.A1(_03482_),
    .A2(_03483_),
    .B1(_03474_),
    .X(_03485_));
 sky130_fd_sc_hd__nand3_1 _09420_ (.A(_03473_),
    .B(_03484_),
    .C(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__and2_1 _09421_ (.A(_03472_),
    .B(_03486_),
    .X(_03488_));
 sky130_fd_sc_hd__nand2_1 _09422_ (.A(_03472_),
    .B(_03486_),
    .Y(_03489_));
 sky130_fd_sc_hd__a21oi_1 _09423_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03435_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21boi_1 _09424_ (.A1(_03482_),
    .A2(_03474_),
    .B1_N(_03483_),
    .Y(_03491_));
 sky130_fd_sc_hd__nand3b_1 _09425_ (.A_N(_02083_),
    .B(_02080_),
    .C(_02077_),
    .Y(_03492_));
 sky130_fd_sc_hd__a21bo_1 _09426_ (.A1(_02077_),
    .A2(_02080_),
    .B1_N(_02083_),
    .X(_03493_));
 sky130_fd_sc_hd__a21boi_1 _09427_ (.A1(_03492_),
    .A2(_03493_),
    .B1_N(_03491_),
    .Y(_03494_));
 sky130_fd_sc_hd__a21bo_1 _09428_ (.A1(_03492_),
    .A2(_03493_),
    .B1_N(_03491_),
    .X(_03495_));
 sky130_fd_sc_hd__a21o_1 _09429_ (.A1(_03484_),
    .A2(_03485_),
    .B1(_03473_),
    .X(_03496_));
 sky130_fd_sc_hd__and3b_1 _09430_ (.A_N(_03491_),
    .B(_03492_),
    .C(_03493_),
    .X(_03497_));
 sky130_fd_sc_hd__nand3b_1 _09431_ (.A_N(_03491_),
    .B(_03492_),
    .C(_03493_),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_03496_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nand3_1 _09433_ (.A(_03495_),
    .B(_03496_),
    .C(_03499_),
    .Y(_03501_));
 sky130_fd_sc_hd__nor4_1 _09434_ (.A(_03489_),
    .B(_03490_),
    .C(_03494_),
    .D(_03500_),
    .Y(_03502_));
 sky130_fd_sc_hd__o2bb2ai_1 _09435_ (.A1_N(_02086_),
    .A2_N(_02087_),
    .B1(_01854_),
    .B2(_02081_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand3_1 _09436_ (.A(_02088_),
    .B(_03503_),
    .C(_03497_),
    .Y(_03504_));
 sky130_fd_sc_hd__o21ai_1 _09437_ (.A1(_03488_),
    .A2(_03501_),
    .B1(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__a21oi_2 _09438_ (.A1(_03434_),
    .A2(_03502_),
    .B1(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__a21oi_2 _09439_ (.A1(_02088_),
    .A2(_03503_),
    .B1(_03497_),
    .Y(_03507_));
 sky130_fd_sc_hd__nor2_2 _09440_ (.A(_03506_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__o2bb2ai_2 _09441_ (.A1_N(_02092_),
    .A2_N(_02089_),
    .B1(_03507_),
    .B2(_03506_),
    .Y(_03510_));
 sky130_fd_sc_hd__o21ai_2 _09442_ (.A1(_02089_),
    .A2(_02092_),
    .B1(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__a31oi_4 _09443_ (.A1(_03510_),
    .A2(_01898_),
    .A3(_02094_),
    .B1(_01896_),
    .Y(_03512_));
 sky130_fd_sc_hd__a22oi_2 _09444_ (.A1(_01690_),
    .A2(_01695_),
    .B1(_01697_),
    .B2(_01699_),
    .Y(_03513_));
 sky130_fd_sc_hd__o21bai_2 _09445_ (.A1(_01698_),
    .A2(_01700_),
    .B1_N(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__o22ai_4 _09446_ (.A1(_01700_),
    .A2(_01698_),
    .B1(_03513_),
    .B2(_03512_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _09447_ (.A(_03515_),
    .B(_01493_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21o_1 _09448_ (.A1(_03515_),
    .A2(_01493_),
    .B1(_01491_),
    .X(_03517_));
 sky130_fd_sc_hd__o211ai_2 _09449_ (.A1(_01126_),
    .A2(_01306_),
    .B1(_01492_),
    .C1(_03516_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand3_2 _09450_ (.A(_03518_),
    .B(_01124_),
    .C(_01308_),
    .Y(_03519_));
 sky130_fd_sc_hd__o41ai_4 _09451_ (.A1(_00933_),
    .A2(_00938_),
    .A3(_01117_),
    .A4(_01121_),
    .B1(_03519_),
    .Y(_03521_));
 sky130_fd_sc_hd__a21bo_1 _09452_ (.A1(_00732_),
    .A2(_00936_),
    .B1_N(_00934_),
    .X(_03522_));
 sky130_fd_sc_hd__a21bo_1 _09453_ (.A1(_00936_),
    .A2(_00937_),
    .B1_N(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__a22oi_4 _09454_ (.A1(_00936_),
    .A2(_00937_),
    .B1(_03521_),
    .B2(_03522_),
    .Y(_03524_));
 sky130_fd_sc_hd__o32ai_4 _09455_ (.A1(_00733_),
    .A2(_00735_),
    .A3(_00736_),
    .B1(_00740_),
    .B2(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand2_1 _09456_ (.A(_00413_),
    .B(_00564_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2b_2 _09457_ (.A_N(_00565_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__a21oi_4 _09458_ (.A1(_03525_),
    .A2(_03526_),
    .B1(_00565_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21bai_4 _09459_ (.A1(_00411_),
    .A2(_03528_),
    .B1_N(_00410_),
    .Y(_03529_));
 sky130_fd_sc_hd__xnor2_2 _09460_ (.A(_00269_),
    .B(_00270_),
    .Y(_03530_));
 sky130_fd_sc_hd__a21oi_4 _09461_ (.A1(_03529_),
    .A2(_03530_),
    .B1(_00271_),
    .Y(_03532_));
 sky130_fd_sc_hd__o21a_1 _09462_ (.A1(_00141_),
    .A2(_03532_),
    .B1(_00139_),
    .X(_03533_));
 sky130_fd_sc_hd__o221ai_4 _09463_ (.A1(_00028_),
    .A2(_00030_),
    .B1(_00141_),
    .B2(_03532_),
    .C1(_00139_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21ai_1 _09464_ (.A1(_00027_),
    .A2(_00029_),
    .B1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__a31oi_4 _09465_ (.A1(_03534_),
    .A2(_05274_),
    .A3(_00031_),
    .B1(_05272_),
    .Y(_03536_));
 sky130_fd_sc_hd__nor2_1 _09466_ (.A(_05098_),
    .B(_05185_),
    .Y(_03537_));
 sky130_fd_sc_hd__or2_2 _09467_ (.A(_05186_),
    .B(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__o21bai_4 _09468_ (.A1(_03538_),
    .A2(_03536_),
    .B1_N(_05186_),
    .Y(_03539_));
 sky130_fd_sc_hd__a21oi_1 _09469_ (.A1(_05012_),
    .A2(_05095_),
    .B1(_05011_),
    .Y(_03540_));
 sky130_fd_sc_hd__a31oi_4 _09470_ (.A1(_03539_),
    .A2(_05096_),
    .A3(_05013_),
    .B1(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__xor2_2 _09471_ (.A(_04805_),
    .B(_04946_),
    .X(_03543_));
 sky130_fd_sc_hd__o32ai_4 _09472_ (.A1(_04719_),
    .A2(_04796_),
    .A3(_04946_),
    .B1(_03543_),
    .B2(_03541_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_2 _09473_ (.A1(_03544_),
    .A2(_04786_),
    .B1(_04758_),
    .Y(_03545_));
 sky130_fd_sc_hd__o21bai_2 _09474_ (.A1(_04180_),
    .A2(_03545_),
    .B1_N(_04158_),
    .Y(_03546_));
 sky130_fd_sc_hd__a21oi_2 _09475_ (.A1(_03546_),
    .A2(_03586_),
    .B1(_03564_),
    .Y(_03547_));
 sky130_fd_sc_hd__o21bai_2 _09476_ (.A1(_03036_),
    .A2(_03547_),
    .B1_N(_03025_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_03548_),
    .B(_02552_),
    .Y(_03549_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_01925_),
    .B(_01947_),
    .Y(_03550_));
 sky130_fd_sc_hd__o211a_1 _09479_ (.A1(_01826_),
    .A2(_01859_),
    .B1(_01881_),
    .C1(_01947_),
    .X(_03551_));
 sky130_fd_sc_hd__o2bb2ai_4 _09480_ (.A1_N(_02519_),
    .A2_N(_03549_),
    .B1(_03550_),
    .B2(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__o211ai_4 _09481_ (.A1(_01914_),
    .A2(_01947_),
    .B1(_01694_),
    .C1(_03552_),
    .Y(_03554_));
 sky130_fd_sc_hd__inv_2 _09482_ (.A(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__a31oi_4 _09483_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_01551_),
    .Y(_03556_));
 sky130_fd_sc_hd__a31o_1 _09484_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_01551_),
    .X(_03557_));
 sky130_fd_sc_hd__xor2_2 _09485_ (.A(_00946_),
    .B(_01001_),
    .X(_03558_));
 sky130_fd_sc_hd__and3b_2 _09486_ (.A_N(_03558_),
    .B(_01089_),
    .C(_01078_),
    .X(_03559_));
 sky130_fd_sc_hd__o2bb2a_1 _09487_ (.A1_N(_01078_),
    .A2_N(_01089_),
    .B1(_00946_),
    .B2(_01012_),
    .X(_03560_));
 sky130_fd_sc_hd__a31o_1 _09488_ (.A1(_00957_),
    .A2(_01001_),
    .A3(_01067_),
    .B1(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__xnor2_2 _09489_ (.A(_01177_),
    .B(_01188_),
    .Y(_03562_));
 sky130_fd_sc_hd__inv_2 _09490_ (.A(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__and3_2 _09491_ (.A(_03559_),
    .B(_01166_),
    .C(_01155_),
    .X(_03565_));
 sky130_fd_sc_hd__nand2_2 _09492_ (.A(_03556_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__xnor2_2 _09493_ (.A(_01199_),
    .B(_01276_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand4b_1 _09494_ (.A_N(_03567_),
    .B(_03554_),
    .C(_01562_),
    .D(_03565_),
    .Y(_03568_));
 sky130_fd_sc_hd__o21ba_1 _09495_ (.A1(_01276_),
    .A2(_01199_),
    .B1_N(_01254_),
    .X(_03569_));
 sky130_fd_sc_hd__xnor2_1 _09496_ (.A(_01353_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__nor2_1 _09497_ (.A(_03567_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand3_2 _09498_ (.A(_03556_),
    .B(_03565_),
    .C(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__o21ai_2 _09499_ (.A1(_01485_),
    .A2(_01496_),
    .B1(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand4_1 _09500_ (.A(_01507_),
    .B(_03556_),
    .C(_03565_),
    .D(_03571_),
    .Y(_03574_));
 sky130_fd_sc_hd__nand2_1 _09501_ (.A(_03566_),
    .B(_03567_),
    .Y(_03576_));
 sky130_fd_sc_hd__nand4_2 _09502_ (.A(_03552_),
    .B(_01694_),
    .C(_01551_),
    .D(_01958_),
    .Y(_03577_));
 sky130_fd_sc_hd__a31o_1 _09503_ (.A1(net21),
    .A2(net53),
    .A3(_01463_),
    .B1(_01485_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2_1 _09504_ (.A(net22),
    .B(net54),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_2 _09505_ (.A(_00297_),
    .B(net24),
    .Y(_03580_));
 sky130_fd_sc_hd__nand2b_2 _09506_ (.A_N(net24),
    .B(net56),
    .Y(_03581_));
 sky130_fd_sc_hd__nand2_2 _09507_ (.A(_03580_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__xnor2_1 _09508_ (.A(_03579_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__nor2_1 _09509_ (.A(_03578_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__and2_1 _09510_ (.A(_03578_),
    .B(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__or2_1 _09511_ (.A(_03584_),
    .B(_03585_),
    .X(_03587_));
 sky130_fd_sc_hd__o211a_1 _09512_ (.A1(_03584_),
    .A2(_03585_),
    .B1(_03559_),
    .C1(_03577_),
    .X(_03588_));
 sky130_fd_sc_hd__nand3_1 _09513_ (.A(_03577_),
    .B(_03587_),
    .C(_03559_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand3b_1 _09514_ (.A_N(_03558_),
    .B(_03554_),
    .C(_01562_),
    .Y(_03590_));
 sky130_fd_sc_hd__a31o_1 _09515_ (.A1(_01562_),
    .A2(_03554_),
    .A3(_03559_),
    .B1(_03562_),
    .X(_03591_));
 sky130_fd_sc_hd__nor4_2 _09516_ (.A(_03563_),
    .B(_03567_),
    .C(_03556_),
    .D(_03589_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand4b_2 _09517_ (.A_N(_03567_),
    .B(_03557_),
    .C(_03562_),
    .D(_03588_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_2 _09518_ (.A(_03568_),
    .B(_03570_),
    .Y(_03594_));
 sky130_fd_sc_hd__o211a_1 _09519_ (.A1(_01364_),
    .A2(_03566_),
    .B1(_03594_),
    .C1(_03592_),
    .X(_03595_));
 sky130_fd_sc_hd__o211ai_2 _09520_ (.A1(_01364_),
    .A2(_03566_),
    .B1(_01507_),
    .C1(_03594_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand4_4 _09521_ (.A(_03592_),
    .B(_03594_),
    .C(_03572_),
    .D(_03573_),
    .Y(_03598_));
 sky130_fd_sc_hd__a2bb2o_2 _09522_ (.A1_N(_00605_),
    .A2_N(_00792_),
    .B1(_00869_),
    .B2(_00737_),
    .X(_03599_));
 sky130_fd_sc_hd__inv_2 _09523_ (.A(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(_00803_),
    .B(_00891_),
    .X(_03601_));
 sky130_fd_sc_hd__nand2_1 _09525_ (.A(_00803_),
    .B(_00891_),
    .Y(_03602_));
 sky130_fd_sc_hd__nor2_4 _09526_ (.A(_00935_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__inv_2 _09527_ (.A(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__or4_1 _09528_ (.A(_05339_),
    .B(_00924_),
    .C(_03599_),
    .D(_03602_),
    .X(_03605_));
 sky130_fd_sc_hd__o21bai_4 _09529_ (.A1(_03593_),
    .A2(_03596_),
    .B1_N(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__xor2_2 _09530_ (.A(_02089_),
    .B(_02092_),
    .X(_03607_));
 sky130_fd_sc_hd__xnor2_4 _09531_ (.A(_03508_),
    .B(_03607_),
    .Y(_03609_));
 sky130_fd_sc_hd__nor2_1 _09532_ (.A(net24),
    .B(net56),
    .Y(_03610_));
 sky130_fd_sc_hd__a2111oi_4 _09533_ (.A1(net22),
    .A2(net54),
    .B1(net56),
    .C1(net24),
    .D1(_03578_),
    .Y(_03611_));
 sky130_fd_sc_hd__or4b_4 _09534_ (.A(net24),
    .B(net56),
    .C(_03578_),
    .D_N(_03579_),
    .X(_03612_));
 sky130_fd_sc_hd__xor2_4 _09535_ (.A(_01898_),
    .B(_03511_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _09536_ (.A0(_03609_),
    .A1(_03613_),
    .S(_03554_),
    .X(_03614_));
 sky130_fd_sc_hd__and2b_4 _09537_ (.A_N(net57),
    .B(net25),
    .X(_03615_));
 sky130_fd_sc_hd__and2b_4 _09538_ (.A_N(net25),
    .B(net57),
    .X(_03616_));
 sky130_fd_sc_hd__or2_4 _09539_ (.A(_03615_),
    .B(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__nor2_8 _09540_ (.A(_03615_),
    .B(_03616_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2b_1 _09541_ (.A_N(net48),
    .B(net16),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_2 _09542_ (.A(_00000_),
    .B(net48),
    .Y(_03621_));
 sky130_fd_sc_hd__o21ai_4 _09543_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_01012_),
    .Y(_03622_));
 sky130_fd_sc_hd__and4b_2 _09544_ (.A_N(_01067_),
    .B(_01133_),
    .C(_01562_),
    .D(_01012_),
    .X(_03623_));
 sky130_fd_sc_hd__nand4b_4 _09545_ (.A_N(_01067_),
    .B(_01562_),
    .C(_01133_),
    .D(_01012_),
    .Y(_03624_));
 sky130_fd_sc_hd__nor2_1 _09546_ (.A(_00968_),
    .B(_03620_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand3_2 _09547_ (.A(_00990_),
    .B(_01034_),
    .C(_01056_),
    .Y(_03626_));
 sky130_fd_sc_hd__o2111a_2 _09548_ (.A1(_00968_),
    .A2(_03620_),
    .B1(_01056_),
    .C1(_01034_),
    .D1(_00990_),
    .X(_03627_));
 sky130_fd_sc_hd__o21ai_2 _09549_ (.A1(net18),
    .A2(_00275_),
    .B1(_01111_),
    .Y(_03628_));
 sky130_fd_sc_hd__o21bai_4 _09550_ (.A1(_03626_),
    .A2(_03625_),
    .B1_N(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__o21ai_2 _09551_ (.A1(_00011_),
    .A2(net51),
    .B1(_03629_),
    .Y(_03631_));
 sky130_fd_sc_hd__o211a_2 _09552_ (.A1(_00011_),
    .A2(net51),
    .B1(_03624_),
    .C1(_03629_),
    .X(_03632_));
 sky130_fd_sc_hd__o211ai_4 _09553_ (.A1(_00011_),
    .A2(net51),
    .B1(_03624_),
    .C1(_03629_),
    .Y(_03633_));
 sky130_fd_sc_hd__or2_1 _09554_ (.A(_01408_),
    .B(_03582_),
    .X(_03634_));
 sky130_fd_sc_hd__and4_4 _09555_ (.A(_01419_),
    .B(_01441_),
    .C(_03580_),
    .D(_03581_),
    .X(_03635_));
 sky130_fd_sc_hd__nand4_4 _09556_ (.A(_01419_),
    .B(_01441_),
    .C(_03580_),
    .D(_03581_),
    .Y(_03636_));
 sky130_fd_sc_hd__o22a_4 _09557_ (.A1(_01210_),
    .A2(_01221_),
    .B1(_01287_),
    .B2(_01309_),
    .X(_03637_));
 sky130_fd_sc_hd__inv_2 _09558_ (.A(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__a211oi_4 _09559_ (.A1(_01298_),
    .A2(_01320_),
    .B1(_01232_),
    .C1(_03636_),
    .Y(_03639_));
 sky130_fd_sc_hd__nand2_4 _09560_ (.A(_03635_),
    .B(_03637_),
    .Y(_03640_));
 sky130_fd_sc_hd__a31oi_4 _09561_ (.A1(_01122_),
    .A2(_03624_),
    .A3(_03629_),
    .B1(_03640_),
    .Y(_03642_));
 sky130_fd_sc_hd__nand2_8 _09562_ (.A(_03633_),
    .B(_03639_),
    .Y(_03643_));
 sky130_fd_sc_hd__nor2_4 _09563_ (.A(net21),
    .B(_00286_),
    .Y(_03644_));
 sky130_fd_sc_hd__and2b_1 _09564_ (.A_N(net52),
    .B(net20),
    .X(_03645_));
 sky130_fd_sc_hd__a21oi_4 _09565_ (.A1(net21),
    .A2(_00286_),
    .B1(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__nor2_1 _09566_ (.A(_03644_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__a21boi_2 _09567_ (.A1(_01430_),
    .A2(_03581_),
    .B1_N(_03580_),
    .Y(_03648_));
 sky130_fd_sc_hd__o31a_4 _09568_ (.A1(_03644_),
    .A2(_03646_),
    .A3(_03636_),
    .B1(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__o31ai_4 _09569_ (.A1(_03644_),
    .A2(_03646_),
    .A3(_03636_),
    .B1(_03648_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21oi_4 _09570_ (.A1(_03633_),
    .A2(_03639_),
    .B1(net115),
    .Y(_03651_));
 sky130_fd_sc_hd__a21o_4 _09571_ (.A1(_03633_),
    .A2(_03639_),
    .B1(net115),
    .X(_03653_));
 sky130_fd_sc_hd__a31o_1 _09572_ (.A1(_01122_),
    .A2(_03624_),
    .A3(_03629_),
    .B1(_01232_),
    .X(_03654_));
 sky130_fd_sc_hd__o2111ai_4 _09573_ (.A1(_00011_),
    .A2(net51),
    .B1(_01232_),
    .C1(_03624_),
    .D1(_03629_),
    .Y(_03655_));
 sky130_fd_sc_hd__a211o_2 _09574_ (.A1(_03654_),
    .A2(_03655_),
    .B1(_03623_),
    .C1(_03653_),
    .X(_03656_));
 sky130_fd_sc_hd__o211ai_4 _09575_ (.A1(_03623_),
    .A2(_03653_),
    .B1(_03654_),
    .C1(_03655_),
    .Y(_03657_));
 sky130_fd_sc_hd__and2_4 _09576_ (.A(_03656_),
    .B(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__nand2_2 _09577_ (.A(_03656_),
    .B(_03657_),
    .Y(_03659_));
 sky130_fd_sc_hd__a21boi_1 _09578_ (.A1(_00979_),
    .A2(_03621_),
    .B1_N(_00990_),
    .Y(_03660_));
 sky130_fd_sc_hd__or3_4 _09579_ (.A(_01023_),
    .B(_01045_),
    .C(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__o211a_1 _09580_ (.A1(net113),
    .A2(net111),
    .B1(_01056_),
    .C1(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__o211ai_4 _09581_ (.A1(net113),
    .A2(net111),
    .B1(_01056_),
    .C1(_03661_),
    .Y(_03664_));
 sky130_fd_sc_hd__o221a_2 _09582_ (.A1(net18),
    .A2(_00275_),
    .B1(_03625_),
    .B2(_03626_),
    .C1(_03651_),
    .X(_03665_));
 sky130_fd_sc_hd__o21a_4 _09583_ (.A1(_03662_),
    .A2(_03665_),
    .B1(_01133_),
    .X(_03666_));
 sky130_fd_sc_hd__o21ai_4 _09584_ (.A1(_03662_),
    .A2(_03665_),
    .B1(_01133_),
    .Y(_03667_));
 sky130_fd_sc_hd__o311a_4 _09585_ (.A1(_01023_),
    .A2(_03627_),
    .A3(_03653_),
    .B1(_03664_),
    .C1(_01144_),
    .X(_03668_));
 sky130_fd_sc_hd__o311ai_4 _09586_ (.A1(_01023_),
    .A2(_03627_),
    .A3(_03653_),
    .B1(_03664_),
    .C1(_01144_),
    .Y(_03669_));
 sky130_fd_sc_hd__o21ai_1 _09587_ (.A1(_03662_),
    .A2(_03665_),
    .B1(_01144_),
    .Y(_03670_));
 sky130_fd_sc_hd__a31o_1 _09588_ (.A1(_01056_),
    .A2(_03653_),
    .A3(_03661_),
    .B1(_01144_),
    .X(_03671_));
 sky130_fd_sc_hd__o21ai_4 _09589_ (.A1(_03665_),
    .A2(_03671_),
    .B1(_03670_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_8 _09590_ (.A(_03667_),
    .B(_03669_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2b_1 _09591_ (.A_N(net20),
    .B(net52),
    .Y(_03675_));
 sky130_fd_sc_hd__a21oi_2 _09592_ (.A1(_03631_),
    .A2(_03675_),
    .B1(_03645_),
    .Y(_03676_));
 sky130_fd_sc_hd__a211o_1 _09593_ (.A1(_01243_),
    .A2(_03633_),
    .B1(_03645_),
    .C1(_03649_),
    .X(_03677_));
 sky130_fd_sc_hd__o21ai_1 _09594_ (.A1(_03676_),
    .A2(_03653_),
    .B1(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_4 _09595_ (.A1(_01287_),
    .A2(_01309_),
    .B1(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__o2111ai_4 _09596_ (.A1(_03676_),
    .A2(_03653_),
    .B1(_01320_),
    .C1(_01298_),
    .D1(_03677_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(_03679_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__and2_2 _09598_ (.A(_03679_),
    .B(_03680_),
    .X(_03682_));
 sky130_fd_sc_hd__and3_1 _09599_ (.A(_03672_),
    .B(_03679_),
    .C(_03680_),
    .X(_03683_));
 sky130_fd_sc_hd__and3_4 _09600_ (.A(_03658_),
    .B(_03679_),
    .C(_03680_),
    .X(_03684_));
 sky130_fd_sc_hd__nand4_4 _09601_ (.A(_03656_),
    .B(_03657_),
    .C(_03679_),
    .D(_03680_),
    .Y(_03686_));
 sky130_fd_sc_hd__nor2_8 _09602_ (.A(_03673_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__or4_4 _09603_ (.A(_03668_),
    .B(_03659_),
    .C(_03666_),
    .D(_03681_),
    .X(_03688_));
 sky130_fd_sc_hd__o21ai_2 _09604_ (.A1(_01023_),
    .A2(_01045_),
    .B1(_03660_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_03661_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__and3_4 _09606_ (.A(_03622_),
    .B(_03690_),
    .C(_03651_),
    .X(_03691_));
 sky130_fd_sc_hd__a221o_2 _09607_ (.A1(_01012_),
    .A2(_01562_),
    .B1(_03661_),
    .B2(_03689_),
    .C1(_03653_),
    .X(_03692_));
 sky130_fd_sc_hd__a21oi_4 _09608_ (.A1(_03651_),
    .A2(_03622_),
    .B1(_03690_),
    .Y(_03693_));
 sky130_fd_sc_hd__a31o_1 _09609_ (.A1(_03622_),
    .A2(_03643_),
    .A3(_03649_),
    .B1(_03690_),
    .X(_03694_));
 sky130_fd_sc_hd__a22oi_4 _09610_ (.A1(_03661_),
    .A2(_03689_),
    .B1(_03651_),
    .B2(_03622_),
    .Y(_03695_));
 sky130_fd_sc_hd__and4_4 _09611_ (.A(_03651_),
    .B(_03661_),
    .C(_03689_),
    .D(_03622_),
    .X(_03697_));
 sky130_fd_sc_hd__nor2_8 _09612_ (.A(_03691_),
    .B(_03693_),
    .Y(_03698_));
 sky130_fd_sc_hd__nor2_8 _09613_ (.A(_03695_),
    .B(_03697_),
    .Y(_03699_));
 sky130_fd_sc_hd__xor2_4 _09614_ (.A(_01001_),
    .B(_03621_),
    .X(_03700_));
 sky130_fd_sc_hd__xnor2_2 _09615_ (.A(_01001_),
    .B(_03621_),
    .Y(_03701_));
 sky130_fd_sc_hd__and3_4 _09616_ (.A(_01551_),
    .B(_03651_),
    .C(_03700_),
    .X(_03702_));
 sky130_fd_sc_hd__o31a_4 _09617_ (.A1(_01562_),
    .A2(net115),
    .A3(net110),
    .B1(_03701_),
    .X(_03703_));
 sky130_fd_sc_hd__o31a_4 _09618_ (.A1(_01562_),
    .A2(net115),
    .A3(net110),
    .B1(_03700_),
    .X(_03704_));
 sky130_fd_sc_hd__a31o_2 _09619_ (.A1(_03643_),
    .A2(_03649_),
    .A3(_01551_),
    .B1(_03701_),
    .X(_03705_));
 sky130_fd_sc_hd__and3_4 _09620_ (.A(_01551_),
    .B(_03651_),
    .C(_03701_),
    .X(_03706_));
 sky130_fd_sc_hd__or4_4 _09621_ (.A(_01562_),
    .B(net115),
    .C(_03700_),
    .D(net110),
    .X(_03708_));
 sky130_fd_sc_hd__nor2_8 _09622_ (.A(_03702_),
    .B(_03703_),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_8 _09623_ (.A(_03704_),
    .B(_03706_),
    .Y(_03710_));
 sky130_fd_sc_hd__a2bb2oi_1 _09624_ (.A1_N(_03644_),
    .A2_N(_03646_),
    .B1(_03637_),
    .B2(_03633_),
    .Y(_03711_));
 sky130_fd_sc_hd__o2bb2ai_4 _09625_ (.A1_N(_03637_),
    .A2_N(_03633_),
    .B1(_03646_),
    .B2(_03644_),
    .Y(_03712_));
 sky130_fd_sc_hd__a211oi_2 _09626_ (.A1(_03633_),
    .A2(_03637_),
    .B1(_03647_),
    .C1(_03649_),
    .Y(_03713_));
 sky130_fd_sc_hd__o221ai_4 _09627_ (.A1(_03644_),
    .A2(_03646_),
    .B1(_03638_),
    .B2(_03632_),
    .C1(_03650_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21o_1 _09628_ (.A1(_03580_),
    .A2(_03581_),
    .B1(_01419_),
    .X(_03715_));
 sky130_fd_sc_hd__nand2_1 _09629_ (.A(_03634_),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__and2_1 _09630_ (.A(_03634_),
    .B(_03715_),
    .X(_03717_));
 sky130_fd_sc_hd__a31o_1 _09631_ (.A1(_03634_),
    .A2(_03650_),
    .A3(_03715_),
    .B1(_01452_),
    .X(_03719_));
 sky130_fd_sc_hd__a21oi_4 _09632_ (.A1(_03714_),
    .A2(_03716_),
    .B1(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__o21bai_4 _09633_ (.A1(_03717_),
    .A2(_03713_),
    .B1_N(_03719_),
    .Y(_03721_));
 sky130_fd_sc_hd__o21ai_4 _09634_ (.A1(_01463_),
    .A2(_03582_),
    .B1(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__o221a_1 _09635_ (.A1(_00011_),
    .A2(net51),
    .B1(_03628_),
    .B2(_03627_),
    .C1(_03637_),
    .X(_03723_));
 sky130_fd_sc_hd__o221ai_4 _09636_ (.A1(_00011_),
    .A2(net51),
    .B1(_03628_),
    .B2(_03627_),
    .C1(_03637_),
    .Y(_03724_));
 sky130_fd_sc_hd__a21oi_4 _09637_ (.A1(_03712_),
    .A2(_03724_),
    .B1(_01463_),
    .Y(_03725_));
 sky130_fd_sc_hd__o21ai_4 _09638_ (.A1(_03711_),
    .A2(_03723_),
    .B1(_01452_),
    .Y(_03726_));
 sky130_fd_sc_hd__o221ai_4 _09639_ (.A1(_01408_),
    .A2(_01430_),
    .B1(_03631_),
    .B2(_03638_),
    .C1(_03712_),
    .Y(_03727_));
 sky130_fd_sc_hd__a31o_2 _09640_ (.A1(_01463_),
    .A2(_03712_),
    .A3(_03724_),
    .B1(_03653_),
    .X(_03728_));
 sky130_fd_sc_hd__o2111ai_4 _09641_ (.A1(_03632_),
    .A2(_03640_),
    .B1(_03727_),
    .C1(_03649_),
    .D1(_03726_),
    .Y(_03730_));
 sky130_fd_sc_hd__a32oi_4 _09642_ (.A1(_03726_),
    .A2(_03727_),
    .A3(_03651_),
    .B1(_03721_),
    .B2(_03636_),
    .Y(_03731_));
 sky130_fd_sc_hd__o2bb2ai_4 _09643_ (.A1_N(_03636_),
    .A2_N(_03721_),
    .B1(_03725_),
    .B2(_03728_),
    .Y(_03732_));
 sky130_fd_sc_hd__nor2_4 _09644_ (.A(_03624_),
    .B(_03640_),
    .Y(_03733_));
 sky130_fd_sc_hd__a2111o_4 _09645_ (.A1(_01298_),
    .A2(_01320_),
    .B1(_03636_),
    .C1(_01232_),
    .D1(_03624_),
    .X(_03734_));
 sky130_fd_sc_hd__o32a_4 _09646_ (.A1(_03624_),
    .A2(_03636_),
    .A3(_03638_),
    .B1(net115),
    .B2(net110),
    .X(_03735_));
 sky130_fd_sc_hd__a31o_4 _09647_ (.A1(_03623_),
    .A2(_03635_),
    .A3(_03637_),
    .B1(_03651_),
    .X(_03736_));
 sky130_fd_sc_hd__a211oi_4 _09648_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_03733_),
    .C1(net65),
    .Y(_03737_));
 sky130_fd_sc_hd__o221ai_4 _09649_ (.A1(_03624_),
    .A2(_03640_),
    .B1(net113),
    .B2(net110),
    .C1(_05339_),
    .Y(_03738_));
 sky130_fd_sc_hd__o2111ai_4 _09650_ (.A1(net113),
    .A2(net111),
    .B1(net45),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03739_));
 sky130_fd_sc_hd__o21ai_2 _09651_ (.A1(_00253_),
    .A2(_03737_),
    .B1(_03739_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_03738_),
    .B(net14),
    .Y(_03742_));
 sky130_fd_sc_hd__a2111o_1 _09653_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_03733_),
    .C1(net46),
    .D1(net65),
    .X(_03743_));
 sky130_fd_sc_hd__o21ai_1 _09654_ (.A1(_00484_),
    .A2(_03738_),
    .B1(_03742_),
    .Y(_03744_));
 sky130_fd_sc_hd__mux4_2 _09655_ (.A0(net46),
    .A1(net45),
    .A2(net14),
    .A3(net13),
    .S0(_01562_),
    .S1(_03738_),
    .X(_03745_));
 sky130_fd_sc_hd__o2111ai_4 _09656_ (.A1(net113),
    .A2(net110),
    .B1(net47),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03746_));
 sky130_fd_sc_hd__o21ai_4 _09657_ (.A1(_00264_),
    .A2(_03737_),
    .B1(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand4_4 _09658_ (.A(_01562_),
    .B(_03722_),
    .C(_03730_),
    .D(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__o41a_4 _09659_ (.A1(net65),
    .A2(_03733_),
    .A3(_00792_),
    .A4(net109),
    .B1(_00880_),
    .X(_03749_));
 sky130_fd_sc_hd__o2111ai_4 _09660_ (.A1(_03725_),
    .A2(_03728_),
    .B1(_03749_),
    .C1(_01551_),
    .D1(_03722_),
    .Y(_03750_));
 sky130_fd_sc_hd__a31o_1 _09661_ (.A1(_03722_),
    .A2(_03730_),
    .A3(_03749_),
    .B1(_01562_),
    .X(_03752_));
 sky130_fd_sc_hd__o2bb2ai_1 _09662_ (.A1_N(_03747_),
    .A2_N(_03731_),
    .B1(_01529_),
    .B2(_00946_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand2_2 _09663_ (.A(_03748_),
    .B(_03750_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand3_2 _09664_ (.A(_03710_),
    .B(_03748_),
    .C(_03750_),
    .Y(_03755_));
 sky130_fd_sc_hd__a22o_2 _09665_ (.A1(_03705_),
    .A2(_03708_),
    .B1(_03745_),
    .B2(_03731_),
    .X(_03756_));
 sky130_fd_sc_hd__o2111ai_4 _09666_ (.A1(_03709_),
    .A2(_03754_),
    .B1(_03756_),
    .C1(_03698_),
    .D1(_03687_),
    .Y(_03757_));
 sky130_fd_sc_hd__a21oi_1 _09667_ (.A1(_03643_),
    .A2(_03649_),
    .B1(net13),
    .Y(_03758_));
 sky130_fd_sc_hd__a31o_2 _09668_ (.A1(_03643_),
    .A2(_03757_),
    .A3(_03649_),
    .B1(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__o2111ai_4 _09669_ (.A1(net112),
    .A2(net111),
    .B1(net42),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03760_));
 sky130_fd_sc_hd__o21ai_2 _09670_ (.A1(_00231_),
    .A2(_03737_),
    .B1(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__o221ai_4 _09671_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_00231_),
    .B2(_03737_),
    .C1(_03760_),
    .Y(_03763_));
 sky130_fd_sc_hd__a31oi_4 _09672_ (.A1(_05339_),
    .A2(_03653_),
    .A3(_03734_),
    .B1(net11),
    .Y(_03764_));
 sky130_fd_sc_hd__o2111a_1 _09673_ (.A1(net112),
    .A2(net111),
    .B1(_00462_),
    .C1(_05339_),
    .D1(_03734_),
    .X(_03765_));
 sky130_fd_sc_hd__a21oi_1 _09674_ (.A1(_00220_),
    .A2(_03738_),
    .B1(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__o21ai_4 _09675_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_01551_),
    .Y(_03767_));
 sky130_fd_sc_hd__o2111ai_1 _09676_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03722_),
    .C1(_03730_),
    .D1(_03761_),
    .Y(_03768_));
 sky130_fd_sc_hd__o2111ai_1 _09677_ (.A1(_03728_),
    .A2(_03725_),
    .B1(_01551_),
    .C1(_03722_),
    .D1(_03766_),
    .Y(_03769_));
 sky130_fd_sc_hd__o2111ai_1 _09678_ (.A1(_01551_),
    .A2(_03761_),
    .B1(net106),
    .C1(_03710_),
    .D1(_03767_),
    .Y(_03770_));
 sky130_fd_sc_hd__a31o_1 _09679_ (.A1(_05339_),
    .A2(_03653_),
    .A3(_03734_),
    .B1(_00198_),
    .X(_03771_));
 sky130_fd_sc_hd__o211ai_2 _09680_ (.A1(_00451_),
    .A2(_03738_),
    .B1(_01551_),
    .C1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__o2111ai_4 _09681_ (.A1(net112),
    .A2(net111),
    .B1(net40),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03774_));
 sky130_fd_sc_hd__o21ai_2 _09682_ (.A1(_00209_),
    .A2(net107),
    .B1(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__o221ai_4 _09683_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_00209_),
    .B2(_03737_),
    .C1(_03774_),
    .Y(_03776_));
 sky130_fd_sc_hd__o2111ai_1 _09684_ (.A1(_01551_),
    .A2(_03775_),
    .B1(_03772_),
    .C1(net106),
    .D1(_03709_),
    .Y(_03777_));
 sky130_fd_sc_hd__a31o_1 _09685_ (.A1(_03731_),
    .A2(_03772_),
    .A3(_03776_),
    .B1(_03710_),
    .X(_03778_));
 sky130_fd_sc_hd__nand3_1 _09686_ (.A(_03710_),
    .B(_03768_),
    .C(_03769_),
    .Y(_03779_));
 sky130_fd_sc_hd__o211ai_4 _09687_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03778_),
    .C1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand3_1 _09688_ (.A(_03699_),
    .B(_03755_),
    .C(_03756_),
    .Y(_03781_));
 sky130_fd_sc_hd__a22o_1 _09689_ (.A1(_03692_),
    .A2(_03694_),
    .B1(_03755_),
    .B2(_03756_),
    .X(_03782_));
 sky130_fd_sc_hd__a2bb2o_1 _09690_ (.A1_N(_03695_),
    .A2_N(_03697_),
    .B1(_03778_),
    .B2(_03779_),
    .X(_03783_));
 sky130_fd_sc_hd__nand4_1 _09691_ (.A(_03783_),
    .B(net108),
    .C(_03782_),
    .D(_03687_),
    .Y(_03785_));
 sky130_fd_sc_hd__o21ai_2 _09692_ (.A1(_00209_),
    .A2(net109),
    .B1(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__a21oi_1 _09693_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03736_),
    .Y(_03787_));
 sky130_fd_sc_hd__a22oi_4 _09694_ (.A1(net40),
    .A2(_03736_),
    .B1(_03787_),
    .B2(_03687_),
    .Y(_03788_));
 sky130_fd_sc_hd__and4_4 _09695_ (.A(_03731_),
    .B(_03749_),
    .C(_01562_),
    .D(_03701_),
    .X(_03789_));
 sky130_fd_sc_hd__o2111ai_4 _09696_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_01551_),
    .C1(_03730_),
    .D1(_03747_),
    .Y(_03790_));
 sky130_fd_sc_hd__o221ai_4 _09697_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03737_),
    .B2(net14),
    .C1(_03743_),
    .Y(_03791_));
 sky130_fd_sc_hd__o2111ai_4 _09698_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03722_),
    .C1(_03730_),
    .D1(_03744_),
    .Y(_03792_));
 sky130_fd_sc_hd__o21ai_1 _09699_ (.A1(_03732_),
    .A2(_03791_),
    .B1(_03790_),
    .Y(_03793_));
 sky130_fd_sc_hd__a2bb2oi_4 _09700_ (.A1_N(_03704_),
    .A2_N(_03706_),
    .B1(_03790_),
    .B2(_03792_),
    .Y(_03794_));
 sky130_fd_sc_hd__a21o_1 _09701_ (.A1(_03793_),
    .A2(_03709_),
    .B1(_03789_),
    .X(_03796_));
 sky130_fd_sc_hd__o22ai_2 _09702_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03789_),
    .B2(_03794_),
    .Y(_03797_));
 sky130_fd_sc_hd__mux4_2 _09703_ (.A0(net42),
    .A1(net41),
    .A2(net10),
    .A3(net9),
    .S0(_01562_),
    .S1(_03738_),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_03798_),
    .B(net106),
    .Y(_03799_));
 sky130_fd_sc_hd__o2111ai_2 _09705_ (.A1(_00253_),
    .A2(_03737_),
    .B1(_03739_),
    .C1(_00957_),
    .D1(_01540_),
    .Y(_03800_));
 sky130_fd_sc_hd__o21ai_2 _09706_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_01562_),
    .Y(_03801_));
 sky130_fd_sc_hd__o2111ai_1 _09707_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_03730_),
    .C1(_01562_),
    .D1(_03766_),
    .Y(_03802_));
 sky130_fd_sc_hd__o2111ai_1 _09708_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_01551_),
    .C1(_03730_),
    .D1(_03741_),
    .Y(_03803_));
 sky130_fd_sc_hd__o2111ai_4 _09709_ (.A1(_01562_),
    .A2(_03741_),
    .B1(_03731_),
    .C1(_03710_),
    .D1(_03801_),
    .Y(_03804_));
 sky130_fd_sc_hd__o211ai_4 _09710_ (.A1(_03704_),
    .A2(_03706_),
    .B1(_03731_),
    .C1(_03798_),
    .Y(_03805_));
 sky130_fd_sc_hd__o21a_1 _09711_ (.A1(_03710_),
    .A2(_03799_),
    .B1(_03804_),
    .X(_03807_));
 sky130_fd_sc_hd__o211ai_4 _09712_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03804_),
    .C1(_03805_),
    .Y(_03808_));
 sky130_fd_sc_hd__o31a_1 _09713_ (.A1(_03698_),
    .A2(_03789_),
    .A3(_03794_),
    .B1(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__o311a_1 _09714_ (.A1(_03698_),
    .A2(_03789_),
    .A3(_03794_),
    .B1(_03808_),
    .C1(_03672_),
    .X(_03810_));
 sky130_fd_sc_hd__nand4_1 _09715_ (.A(_03809_),
    .B(_03735_),
    .C(_03684_),
    .D(_03672_),
    .Y(_03811_));
 sky130_fd_sc_hd__o21ai_2 _09716_ (.A1(_00451_),
    .A2(_03735_),
    .B1(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__a21oi_1 _09717_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00198_),
    .Y(_03813_));
 sky130_fd_sc_hd__a31o_1 _09718_ (.A1(_03809_),
    .A2(_03687_),
    .A3(net109),
    .B1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__a31oi_1 _09719_ (.A1(_03809_),
    .A2(_03687_),
    .A3(net109),
    .B1(_03813_),
    .Y(_03815_));
 sky130_fd_sc_hd__o211ai_1 _09720_ (.A1(_00451_),
    .A2(_03735_),
    .B1(_03811_),
    .C1(_03814_),
    .Y(_03816_));
 sky130_fd_sc_hd__o2bb2ai_1 _09721_ (.A1_N(_03786_),
    .A2_N(_03788_),
    .B1(_03815_),
    .B2(_03812_),
    .Y(_03818_));
 sky130_fd_sc_hd__nand2_1 _09722_ (.A(_03812_),
    .B(_03815_),
    .Y(_03819_));
 sky130_fd_sc_hd__a31oi_2 _09723_ (.A1(_03801_),
    .A2(_03731_),
    .A3(_03800_),
    .B1(_03710_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand3_2 _09724_ (.A(_03802_),
    .B(_03803_),
    .C(_03709_),
    .Y(_03821_));
 sky130_fd_sc_hd__o211a_1 _09725_ (.A1(_03732_),
    .A2(_03791_),
    .B1(_03790_),
    .C1(_03710_),
    .X(_03822_));
 sky130_fd_sc_hd__o211ai_4 _09726_ (.A1(_03732_),
    .A2(_03791_),
    .B1(_03790_),
    .C1(_03710_),
    .Y(_03823_));
 sky130_fd_sc_hd__o211ai_2 _09727_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03821_),
    .C1(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__o2111ai_4 _09728_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03700_),
    .C1(_03731_),
    .D1(_03749_),
    .Y(_03825_));
 sky130_fd_sc_hd__a21oi_1 _09729_ (.A1(_03692_),
    .A2(_03694_),
    .B1(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__a31oi_2 _09730_ (.A1(_03698_),
    .A2(_03821_),
    .A3(_03823_),
    .B1(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a31o_1 _09731_ (.A1(_03698_),
    .A2(_03821_),
    .A3(_03823_),
    .B1(_03826_),
    .X(_03829_));
 sky130_fd_sc_hd__a21oi_1 _09732_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00462_),
    .Y(_03830_));
 sky130_fd_sc_hd__a31o_1 _09733_ (.A1(_03829_),
    .A2(_03735_),
    .A3(_03687_),
    .B1(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__a31oi_1 _09734_ (.A1(_03829_),
    .A2(_03735_),
    .A3(_03687_),
    .B1(_03830_),
    .Y(_03832_));
 sky130_fd_sc_hd__o21ai_1 _09735_ (.A1(net115),
    .A2(net110),
    .B1(net11),
    .Y(_03833_));
 sky130_fd_sc_hd__o31a_2 _09736_ (.A1(_03653_),
    .A2(_03688_),
    .A3(_03827_),
    .B1(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__a22oi_4 _09737_ (.A1(_03705_),
    .A2(_03708_),
    .B1(_03748_),
    .B2(_03750_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand4_2 _09738_ (.A(_03699_),
    .B(_03753_),
    .C(_03709_),
    .D(_03752_),
    .Y(_03836_));
 sky130_fd_sc_hd__o2111ai_4 _09739_ (.A1(_01551_),
    .A2(_03761_),
    .B1(net106),
    .C1(_03709_),
    .D1(_03767_),
    .Y(_03837_));
 sky130_fd_sc_hd__o211ai_2 _09740_ (.A1(_03702_),
    .A2(_03703_),
    .B1(_03731_),
    .C1(_03745_),
    .Y(_03838_));
 sky130_fd_sc_hd__a21oi_2 _09741_ (.A1(_03745_),
    .A2(_03731_),
    .B1(_03709_),
    .Y(_03840_));
 sky130_fd_sc_hd__a31oi_4 _09742_ (.A1(_03767_),
    .A2(_03731_),
    .A3(_03763_),
    .B1(_03710_),
    .Y(_03841_));
 sky130_fd_sc_hd__o211ai_2 _09743_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03837_),
    .C1(_03838_),
    .Y(_03842_));
 sky130_fd_sc_hd__o31a_2 _09744_ (.A1(_03699_),
    .A2(_03840_),
    .A3(_03841_),
    .B1(_03836_),
    .X(_03843_));
 sky130_fd_sc_hd__o211a_1 _09745_ (.A1(_03698_),
    .A2(_03835_),
    .B1(_03683_),
    .C1(_03842_),
    .X(_03844_));
 sky130_fd_sc_hd__o21ai_2 _09746_ (.A1(net114),
    .A2(net110),
    .B1(net10),
    .Y(_03845_));
 sky130_fd_sc_hd__o31ai_2 _09747_ (.A1(_03653_),
    .A2(_03688_),
    .A3(_03843_),
    .B1(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__o21ai_1 _09748_ (.A1(net109),
    .A2(_03733_),
    .B1(net42),
    .Y(_03847_));
 sky130_fd_sc_hd__o31ai_2 _09749_ (.A1(_03688_),
    .A2(_03736_),
    .A3(_03843_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__o311ai_2 _09750_ (.A1(_03688_),
    .A2(_03736_),
    .A3(_03843_),
    .B1(_03847_),
    .C1(_03846_),
    .Y(_03849_));
 sky130_fd_sc_hd__o21a_1 _09751_ (.A1(_03831_),
    .A2(_03834_),
    .B1(_03849_),
    .X(_03851_));
 sky130_fd_sc_hd__o21ai_1 _09752_ (.A1(net109),
    .A2(_03733_),
    .B1(net45),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_4 _09753_ (.A1(_03736_),
    .A2(_03757_),
    .B1(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _09754_ (.A(_03831_),
    .B(_03834_),
    .Y(_03854_));
 sky130_fd_sc_hd__a22o_1 _09755_ (.A1(_03759_),
    .A2(_03853_),
    .B1(_03834_),
    .B2(_03831_),
    .X(_03855_));
 sky130_fd_sc_hd__a21oi_1 _09756_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00484_),
    .Y(_03856_));
 sky130_fd_sc_hd__a41oi_4 _09757_ (.A1(_03796_),
    .A2(_03735_),
    .A3(_03698_),
    .A4(_03687_),
    .B1(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__a21oi_1 _09758_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00242_),
    .Y(_03858_));
 sky130_fd_sc_hd__a41o_1 _09759_ (.A1(_03796_),
    .A2(_03698_),
    .A3(_03687_),
    .A4(net109),
    .B1(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__nand4_2 _09760_ (.A(_03687_),
    .B(_03698_),
    .C(_03709_),
    .D(_03754_),
    .Y(_03860_));
 sky130_fd_sc_hd__o21ai_1 _09761_ (.A1(net114),
    .A2(net110),
    .B1(net15),
    .Y(_03862_));
 sky130_fd_sc_hd__o21ai_1 _09762_ (.A1(_03653_),
    .A2(_03860_),
    .B1(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__a21oi_1 _09763_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net47),
    .Y(_03864_));
 sky130_fd_sc_hd__a31oi_2 _09764_ (.A1(_03687_),
    .A2(_03698_),
    .A3(_03835_),
    .B1(_03736_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21oi_1 _09765_ (.A1(_03860_),
    .A2(_03735_),
    .B1(_03864_),
    .Y(_03866_));
 sky130_fd_sc_hd__o21ai_1 _09766_ (.A1(_03864_),
    .A2(_03865_),
    .B1(_03863_),
    .Y(_03867_));
 sky130_fd_sc_hd__o211ai_1 _09767_ (.A1(_03653_),
    .A2(_03860_),
    .B1(_03862_),
    .C1(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__o2111a_1 _09768_ (.A1(_03857_),
    .A2(_03859_),
    .B1(_03867_),
    .C1(_03868_),
    .D1(_03733_),
    .X(_03869_));
 sky130_fd_sc_hd__o311ai_2 _09769_ (.A1(_03653_),
    .A2(_03688_),
    .A3(_03843_),
    .B1(_03845_),
    .C1(_03848_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_03859_),
    .B(_03857_),
    .Y(_03871_));
 sky130_fd_sc_hd__a2bb2o_1 _09771_ (.A1_N(_03759_),
    .A2_N(_03853_),
    .B1(_03857_),
    .B2(_03859_),
    .X(_03873_));
 sky130_fd_sc_hd__o2111a_1 _09772_ (.A1(_03759_),
    .A2(_03853_),
    .B1(_03819_),
    .C1(_03816_),
    .D1(_03869_),
    .X(_03874_));
 sky130_fd_sc_hd__o2111a_1 _09773_ (.A1(_03831_),
    .A2(_03834_),
    .B1(_03849_),
    .C1(_03870_),
    .D1(_03871_),
    .X(_03875_));
 sky130_fd_sc_hd__a22oi_1 _09774_ (.A1(_03853_),
    .A2(_03759_),
    .B1(_03786_),
    .B2(_03788_),
    .Y(_03876_));
 sky130_fd_sc_hd__o211a_1 _09775_ (.A1(_03786_),
    .A2(_03788_),
    .B1(_03854_),
    .C1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__nand3_1 _09776_ (.A(_03874_),
    .B(_03875_),
    .C(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21oi_1 _09777_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00176_),
    .Y(_03879_));
 sky130_fd_sc_hd__and3_1 _09778_ (.A(_03692_),
    .B(_03694_),
    .C(_03700_),
    .X(_03880_));
 sky130_fd_sc_hd__o2111ai_4 _09779_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03731_),
    .C1(_03749_),
    .D1(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__a21oi_4 _09780_ (.A1(_03667_),
    .A2(_03669_),
    .B1(_03686_),
    .Y(_03882_));
 sky130_fd_sc_hd__or3_1 _09781_ (.A(_03681_),
    .B(_03659_),
    .C(_03672_),
    .X(_03884_));
 sky130_fd_sc_hd__a211o_1 _09782_ (.A1(_03667_),
    .A2(_03669_),
    .B1(_03686_),
    .C1(_03881_),
    .X(_03885_));
 sky130_fd_sc_hd__o2111ai_4 _09783_ (.A1(_00209_),
    .A2(net107),
    .B1(_03774_),
    .C1(_00957_),
    .D1(_01540_),
    .Y(_03886_));
 sky130_fd_sc_hd__o2111ai_4 _09784_ (.A1(net112),
    .A2(net111),
    .B1(net39),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03887_));
 sky130_fd_sc_hd__o21ai_1 _09785_ (.A1(_00176_),
    .A2(net107),
    .B1(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__o221ai_4 _09786_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_00176_),
    .B2(net107),
    .C1(_03887_),
    .Y(_03889_));
 sky130_fd_sc_hd__o2111ai_1 _09787_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_03730_),
    .C1(_03888_),
    .D1(_01562_),
    .Y(_03890_));
 sky130_fd_sc_hd__o2111ai_1 _09788_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_01551_),
    .C1(_03730_),
    .D1(_03775_),
    .Y(_03891_));
 sky130_fd_sc_hd__o2111ai_2 _09789_ (.A1(_01562_),
    .A2(_03775_),
    .B1(net106),
    .C1(_03889_),
    .D1(_03709_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand3_1 _09790_ (.A(_03890_),
    .B(_03891_),
    .C(_03709_),
    .Y(_03893_));
 sky130_fd_sc_hd__o2bb2ai_1 _09791_ (.A1_N(net106),
    .A2_N(_03798_),
    .B1(_03702_),
    .B2(_03703_),
    .Y(_03895_));
 sky130_fd_sc_hd__o21ai_2 _09792_ (.A1(_03709_),
    .A2(_03799_),
    .B1(_03892_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand3_1 _09793_ (.A(_03893_),
    .B(_03895_),
    .C(_03698_),
    .Y(_03897_));
 sky130_fd_sc_hd__o211ai_1 _09794_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03821_),
    .C1(_03823_),
    .Y(_03898_));
 sky130_fd_sc_hd__o22ai_4 _09795_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03820_),
    .B2(_03822_),
    .Y(_03899_));
 sky130_fd_sc_hd__o211ai_1 _09796_ (.A1(_03709_),
    .A2(_03799_),
    .B1(_03892_),
    .C1(_03698_),
    .Y(_03900_));
 sky130_fd_sc_hd__nand3_1 _09797_ (.A(_03899_),
    .B(_03900_),
    .C(_03687_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand3_2 _09798_ (.A(_03898_),
    .B(_03672_),
    .C(_03897_),
    .Y(_03902_));
 sky130_fd_sc_hd__a21oi_2 _09799_ (.A1(_03673_),
    .A2(_03881_),
    .B1(_03686_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_1 _09800_ (.A1(net114),
    .A2(net110),
    .B1(_00176_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand3_1 _09801_ (.A(_03901_),
    .B(net108),
    .C(_03885_),
    .Y(_03906_));
 sky130_fd_sc_hd__a31oi_2 _09802_ (.A1(_03902_),
    .A2(_03903_),
    .A3(net109),
    .B1(_03879_),
    .Y(_03907_));
 sky130_fd_sc_hd__a31o_1 _09803_ (.A1(_03902_),
    .A2(_03903_),
    .A3(net109),
    .B1(_03879_),
    .X(_03908_));
 sky130_fd_sc_hd__a21oi_1 _09804_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00440_),
    .Y(_03909_));
 sky130_fd_sc_hd__a31oi_1 _09805_ (.A1(_03902_),
    .A2(_03903_),
    .A3(_03735_),
    .B1(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__a31o_1 _09806_ (.A1(_03902_),
    .A2(_03903_),
    .A3(_03735_),
    .B1(_03909_),
    .X(_03911_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(_03911_),
    .B(_03907_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand4_2 _09808_ (.A(_03754_),
    .B(_03882_),
    .C(_03698_),
    .D(_03709_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand4_2 _09809_ (.A(net106),
    .B(_03772_),
    .C(_03776_),
    .D(_03710_),
    .Y(_03914_));
 sky130_fd_sc_hd__o211ai_2 _09810_ (.A1(_00176_),
    .A2(net107),
    .B1(_03887_),
    .C1(_01551_),
    .Y(_03915_));
 sky130_fd_sc_hd__o2111ai_2 _09811_ (.A1(net112),
    .A2(net111),
    .B1(net38),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03917_));
 sky130_fd_sc_hd__o221ai_4 _09812_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_00187_),
    .B2(net107),
    .C1(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__nand4_2 _09813_ (.A(_03709_),
    .B(net106),
    .C(_03915_),
    .D(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__o211ai_2 _09814_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03837_),
    .C1(_03838_),
    .Y(_03920_));
 sky130_fd_sc_hd__o211ai_2 _09815_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03914_),
    .C1(_03919_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand4_2 _09816_ (.A(_03920_),
    .B(_03921_),
    .C(_03672_),
    .D(_03684_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21oi_1 _09817_ (.A1(_03643_),
    .A2(_03649_),
    .B1(net6),
    .Y(_03923_));
 sky130_fd_sc_hd__a31o_1 _09818_ (.A1(_03922_),
    .A2(net109),
    .A3(_03913_),
    .B1(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__a31oi_1 _09819_ (.A1(_03922_),
    .A2(net109),
    .A3(_03913_),
    .B1(_03923_),
    .Y(_03925_));
 sky130_fd_sc_hd__a21oi_1 _09820_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net38),
    .Y(_03926_));
 sky130_fd_sc_hd__a31o_1 _09821_ (.A1(_03922_),
    .A2(_03735_),
    .A3(_03913_),
    .B1(_03926_),
    .X(_03928_));
 sky130_fd_sc_hd__a31oi_1 _09822_ (.A1(_03922_),
    .A2(_03735_),
    .A3(_03913_),
    .B1(_03926_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _09823_ (.A(_03928_),
    .B(_03925_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_03924_),
    .B(_03929_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand3_1 _09825_ (.A(_03910_),
    .B(_03906_),
    .C(_03904_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand4_2 _09826_ (.A(_03912_),
    .B(_03930_),
    .C(_03931_),
    .D(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand4_2 _09827_ (.A(_03755_),
    .B(_03882_),
    .C(_03756_),
    .D(_03698_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand4_1 _09828_ (.A(net106),
    .B(_03915_),
    .C(_03918_),
    .D(_03710_),
    .Y(_03935_));
 sky130_fd_sc_hd__a31oi_1 _09829_ (.A1(_05339_),
    .A2(_03653_),
    .A3(_03734_),
    .B1(_00165_),
    .Y(_03936_));
 sky130_fd_sc_hd__o2111a_1 _09830_ (.A1(net112),
    .A2(net111),
    .B1(net36),
    .C1(_05339_),
    .D1(_03734_),
    .X(_03937_));
 sky130_fd_sc_hd__a21oi_1 _09831_ (.A1(net4),
    .A2(_03738_),
    .B1(_03937_),
    .Y(_03939_));
 sky130_fd_sc_hd__mux4_2 _09832_ (.A0(net37),
    .A1(net36),
    .A2(net5),
    .A3(net4),
    .S0(_01562_),
    .S1(_03738_),
    .X(_03940_));
 sky130_fd_sc_hd__o211ai_1 _09833_ (.A1(_03704_),
    .A2(_03706_),
    .B1(net106),
    .C1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__o2bb2ai_1 _09834_ (.A1_N(net106),
    .A2_N(_03940_),
    .B1(_03704_),
    .B2(_03706_),
    .Y(_03942_));
 sky130_fd_sc_hd__a31o_1 _09835_ (.A1(net106),
    .A2(_03915_),
    .A3(_03918_),
    .B1(_03709_),
    .X(_03943_));
 sky130_fd_sc_hd__o211ai_2 _09836_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03770_),
    .C1(_03777_),
    .Y(_03944_));
 sky130_fd_sc_hd__o211ai_2 _09837_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03935_),
    .C1(_03941_),
    .Y(_03945_));
 sky130_fd_sc_hd__nand4_2 _09838_ (.A(_03944_),
    .B(_03945_),
    .C(_03672_),
    .D(_03684_),
    .Y(_03946_));
 sky130_fd_sc_hd__a21oi_1 _09839_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net36),
    .Y(_03947_));
 sky130_fd_sc_hd__a31oi_1 _09840_ (.A1(_03946_),
    .A2(_03735_),
    .A3(_03934_),
    .B1(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a31o_1 _09841_ (.A1(_03946_),
    .A2(_03735_),
    .A3(_03934_),
    .B1(_03947_),
    .X(_03950_));
 sky130_fd_sc_hd__nand3_1 _09842_ (.A(_03946_),
    .B(net109),
    .C(_03934_),
    .Y(_03951_));
 sky130_fd_sc_hd__o21ai_2 _09843_ (.A1(net4),
    .A2(net109),
    .B1(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand2_1 _09844_ (.A(_03948_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__o211ai_1 _09845_ (.A1(net4),
    .A2(net109),
    .B1(_03950_),
    .C1(_03951_),
    .Y(_03954_));
 sky130_fd_sc_hd__o211ai_4 _09846_ (.A1(_03789_),
    .A2(_03794_),
    .B1(_03882_),
    .C1(_03698_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand4_4 _09847_ (.A(net106),
    .B(_03886_),
    .C(_03889_),
    .D(_03710_),
    .Y(_03956_));
 sky130_fd_sc_hd__mux4_2 _09848_ (.A0(net38),
    .A1(net37),
    .A2(net6),
    .A3(net5),
    .S0(_01562_),
    .S1(_03738_),
    .X(_03957_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_03957_),
    .B(net106),
    .Y(_03958_));
 sky130_fd_sc_hd__o211ai_2 _09850_ (.A1(_03704_),
    .A2(_03706_),
    .B1(net106),
    .C1(_03957_),
    .Y(_03959_));
 sky130_fd_sc_hd__o211ai_4 _09851_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03804_),
    .C1(_03805_),
    .Y(_03961_));
 sky130_fd_sc_hd__o211ai_4 _09852_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03956_),
    .C1(_03959_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand4_4 _09853_ (.A(_03961_),
    .B(_03962_),
    .C(_03672_),
    .D(_03684_),
    .Y(_03963_));
 sky130_fd_sc_hd__a21oi_1 _09854_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net37),
    .Y(_03964_));
 sky130_fd_sc_hd__a31o_1 _09855_ (.A1(_03955_),
    .A2(_03963_),
    .A3(_03735_),
    .B1(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a31oi_1 _09856_ (.A1(_03955_),
    .A2(_03963_),
    .A3(_03735_),
    .B1(_03964_),
    .Y(_03966_));
 sky130_fd_sc_hd__a21oi_1 _09857_ (.A1(_03643_),
    .A2(_03649_),
    .B1(net5),
    .Y(_03967_));
 sky130_fd_sc_hd__a31o_1 _09858_ (.A1(_03955_),
    .A2(_03963_),
    .A3(net109),
    .B1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__a31oi_2 _09859_ (.A1(_03955_),
    .A2(_03963_),
    .A3(net109),
    .B1(_03967_),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_03965_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _09861_ (.A(_03968_),
    .B(_03966_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand4_1 _09862_ (.A(_03953_),
    .B(_03954_),
    .C(_03970_),
    .D(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__o211ai_1 _09863_ (.A1(_03965_),
    .A2(_03969_),
    .B1(_03953_),
    .C1(_03954_),
    .Y(_03974_));
 sky130_fd_sc_hd__nor2_1 _09864_ (.A(_03933_),
    .B(_03973_),
    .Y(_03975_));
 sky130_fd_sc_hd__a211o_1 _09865_ (.A1(_03965_),
    .A2(_03969_),
    .B1(_03974_),
    .C1(_03933_),
    .X(_03976_));
 sky130_fd_sc_hd__o211ai_1 _09866_ (.A1(_03702_),
    .A2(_03703_),
    .B1(net106),
    .C1(_03940_),
    .Y(_03977_));
 sky130_fd_sc_hd__o2111ai_1 _09867_ (.A1(net112),
    .A2(net111),
    .B1(net35),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03978_));
 sky130_fd_sc_hd__o21a_1 _09868_ (.A1(_00132_),
    .A2(net107),
    .B1(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__o21ai_1 _09869_ (.A1(_00132_),
    .A2(net107),
    .B1(_03978_),
    .Y(_03980_));
 sky130_fd_sc_hd__o2111ai_1 _09870_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_01551_),
    .C1(_03730_),
    .D1(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__o2111ai_2 _09871_ (.A1(net112),
    .A2(net111),
    .B1(net34),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_03983_));
 sky130_fd_sc_hd__a21boi_1 _09872_ (.A1(net2),
    .A2(_03738_),
    .B1_N(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__o21ai_2 _09873_ (.A1(_00143_),
    .A2(net107),
    .B1(_03983_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand4_1 _09874_ (.A(_01562_),
    .B(_03722_),
    .C(_03730_),
    .D(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__o22ai_1 _09875_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03984_),
    .B2(_03732_),
    .Y(_03987_));
 sky130_fd_sc_hd__o21ai_1 _09876_ (.A1(_03979_),
    .A2(_03732_),
    .B1(_01551_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand3_1 _09877_ (.A(_03988_),
    .B(_03709_),
    .C(_03987_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand3_1 _09878_ (.A(_03986_),
    .B(_03709_),
    .C(_03981_),
    .Y(_03990_));
 sky130_fd_sc_hd__o2bb2ai_1 _09879_ (.A1_N(net106),
    .A2_N(_03940_),
    .B1(_03702_),
    .B2(_03703_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand3_1 _09880_ (.A(_03990_),
    .B(_03991_),
    .C(_03698_),
    .Y(_03992_));
 sky130_fd_sc_hd__a22o_1 _09881_ (.A1(_03692_),
    .A2(_03694_),
    .B1(_03914_),
    .B2(_03919_),
    .X(_03994_));
 sky130_fd_sc_hd__nand3_1 _09882_ (.A(_03699_),
    .B(_03914_),
    .C(_03919_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand3_1 _09883_ (.A(_03989_),
    .B(_03698_),
    .C(_03977_),
    .Y(_03996_));
 sky130_fd_sc_hd__nand3_1 _09884_ (.A(_03996_),
    .B(_03687_),
    .C(_03995_),
    .Y(_03997_));
 sky130_fd_sc_hd__o2111ai_1 _09885_ (.A1(_03698_),
    .A2(_03835_),
    .B1(_03842_),
    .C1(_03684_),
    .D1(_03673_),
    .Y(_03998_));
 sky130_fd_sc_hd__o311ai_4 _09886_ (.A1(_03699_),
    .A2(_03840_),
    .A3(_03841_),
    .B1(_03836_),
    .C1(_03673_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand3_1 _09887_ (.A(_03994_),
    .B(_03672_),
    .C(_03992_),
    .Y(_04000_));
 sky130_fd_sc_hd__a21oi_1 _09888_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00143_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand3_1 _09889_ (.A(_03997_),
    .B(_03998_),
    .C(net108),
    .Y(_04002_));
 sky130_fd_sc_hd__a41oi_1 _09890_ (.A1(_03999_),
    .A2(_04000_),
    .A3(net108),
    .A4(_03684_),
    .B1(_04001_),
    .Y(_04003_));
 sky130_fd_sc_hd__a41o_1 _09891_ (.A1(_03999_),
    .A2(_04000_),
    .A3(net108),
    .A4(_03684_),
    .B1(_04001_),
    .X(_04005_));
 sky130_fd_sc_hd__o211ai_1 _09892_ (.A1(_03884_),
    .A2(_03843_),
    .B1(_03735_),
    .C1(_03997_),
    .Y(_04006_));
 sky130_fd_sc_hd__o21ai_1 _09893_ (.A1(net108),
    .A2(_03733_),
    .B1(_00418_),
    .Y(_04007_));
 sky130_fd_sc_hd__a21oi_1 _09894_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00418_),
    .Y(_04008_));
 sky130_fd_sc_hd__nand4_1 _09895_ (.A(_03999_),
    .B(_04000_),
    .C(_03684_),
    .D(_03735_),
    .Y(_04009_));
 sky130_fd_sc_hd__a41o_1 _09896_ (.A1(_03999_),
    .A2(_04000_),
    .A3(_03684_),
    .A4(_03735_),
    .B1(_04008_),
    .X(_04010_));
 sky130_fd_sc_hd__o21ai_1 _09897_ (.A1(net34),
    .A2(_03735_),
    .B1(_04006_),
    .Y(_04011_));
 sky130_fd_sc_hd__o211ai_1 _09898_ (.A1(net2),
    .A2(net108),
    .B1(_04002_),
    .C1(_04009_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand3_1 _09899_ (.A(_04003_),
    .B(_04006_),
    .C(_04007_),
    .Y(_04013_));
 sky130_fd_sc_hd__a21oi_1 _09900_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00132_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand3_1 _09901_ (.A(_03699_),
    .B(_03893_),
    .C(_03895_),
    .Y(_04016_));
 sky130_fd_sc_hd__o21ai_1 _09902_ (.A1(_03936_),
    .A2(_03937_),
    .B1(_01551_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand4_1 _09903_ (.A(_01562_),
    .B(_03722_),
    .C(_03730_),
    .D(_03980_),
    .Y(_04018_));
 sky130_fd_sc_hd__o22ai_2 _09904_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03979_),
    .B2(_03732_),
    .Y(_04019_));
 sky130_fd_sc_hd__o21ai_1 _09905_ (.A1(_03939_),
    .A2(_03732_),
    .B1(_01551_),
    .Y(_04020_));
 sky130_fd_sc_hd__o211ai_2 _09906_ (.A1(_03704_),
    .A2(_03706_),
    .B1(_04019_),
    .C1(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__o211ai_1 _09907_ (.A1(_03732_),
    .A2(_04017_),
    .B1(_04018_),
    .C1(_03709_),
    .Y(_04022_));
 sky130_fd_sc_hd__a2bb2o_1 _09908_ (.A1_N(_03702_),
    .A2_N(_03703_),
    .B1(net106),
    .B2(_03957_),
    .X(_04023_));
 sky130_fd_sc_hd__nand3_1 _09909_ (.A(_04022_),
    .B(_04023_),
    .C(_03698_),
    .Y(_04024_));
 sky130_fd_sc_hd__o211ai_1 _09910_ (.A1(_03709_),
    .A2(_03958_),
    .B1(_03698_),
    .C1(_04021_),
    .Y(_04025_));
 sky130_fd_sc_hd__o2111ai_1 _09911_ (.A1(_03698_),
    .A2(_03896_),
    .B1(_03672_),
    .C1(_03684_),
    .D1(_04025_),
    .Y(_04027_));
 sky130_fd_sc_hd__o211ai_4 _09912_ (.A1(_03825_),
    .A2(_03698_),
    .B1(_03673_),
    .C1(_03824_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand3_2 _09913_ (.A(_04024_),
    .B(_03672_),
    .C(_04016_),
    .Y(_04029_));
 sky130_fd_sc_hd__a41oi_2 _09914_ (.A1(_04028_),
    .A2(_04029_),
    .A3(net109),
    .A4(_03684_),
    .B1(_04014_),
    .Y(_04030_));
 sky130_fd_sc_hd__a41o_1 _09915_ (.A1(_04029_),
    .A2(net109),
    .A3(_04028_),
    .A4(_03684_),
    .B1(_04014_),
    .X(_04031_));
 sky130_fd_sc_hd__a21oi_1 _09916_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00407_),
    .Y(_04032_));
 sky130_fd_sc_hd__o211ai_1 _09917_ (.A1(_03884_),
    .A2(_03827_),
    .B1(_03735_),
    .C1(_04027_),
    .Y(_04033_));
 sky130_fd_sc_hd__a41oi_4 _09918_ (.A1(_04028_),
    .A2(_04029_),
    .A3(_03684_),
    .A4(_03735_),
    .B1(_04032_),
    .Y(_04034_));
 sky130_fd_sc_hd__o211ai_1 _09919_ (.A1(net35),
    .A2(_03735_),
    .B1(_04033_),
    .C1(_04030_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _09920_ (.A(_04031_),
    .B(_04034_),
    .Y(_04036_));
 sky130_fd_sc_hd__o2111a_1 _09921_ (.A1(_04008_),
    .A2(_04012_),
    .B1(_04013_),
    .C1(_04035_),
    .D1(_04036_),
    .X(_04038_));
 sky130_fd_sc_hd__a21oi_2 _09922_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00121_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _09923_ (.A(_03738_),
    .B(net32),
    .Y(_04040_));
 sky130_fd_sc_hd__o2111ai_1 _09924_ (.A1(net112),
    .A2(net111),
    .B1(net64),
    .C1(_05339_),
    .D1(_03734_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_1 _09925_ (.A1(_00110_),
    .A2(net107),
    .B1(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__mux4_1 _09926_ (.A0(net64),
    .A1(net63),
    .A2(net32),
    .A3(net31),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04043_));
 sky130_fd_sc_hd__a22o_1 _09927_ (.A1(_03705_),
    .A2(_03708_),
    .B1(_04043_),
    .B2(net106),
    .X(_04044_));
 sky130_fd_sc_hd__nand3_1 _09928_ (.A(_03710_),
    .B(_03981_),
    .C(_03986_),
    .Y(_04045_));
 sky130_fd_sc_hd__o211ai_2 _09929_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_04044_),
    .C1(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__o211ai_2 _09930_ (.A1(_03691_),
    .A2(_03693_),
    .B1(_03942_),
    .C1(_03943_),
    .Y(_04047_));
 sky130_fd_sc_hd__o211ai_4 _09931_ (.A1(_03666_),
    .A2(_03668_),
    .B1(_03780_),
    .C1(_03781_),
    .Y(_04049_));
 sky130_fd_sc_hd__nand3_1 _09932_ (.A(_04046_),
    .B(_04047_),
    .C(_03672_),
    .Y(_04050_));
 sky130_fd_sc_hd__a41oi_2 _09933_ (.A1(_04049_),
    .A2(_04050_),
    .A3(net108),
    .A4(_03684_),
    .B1(_04039_),
    .Y(_04051_));
 sky130_fd_sc_hd__a41o_1 _09934_ (.A1(_04049_),
    .A2(_04050_),
    .A3(net108),
    .A4(_03684_),
    .B1(_04039_),
    .X(_04052_));
 sky130_fd_sc_hd__a21oi_1 _09935_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00396_),
    .Y(_04053_));
 sky130_fd_sc_hd__a41o_1 _09936_ (.A1(_04049_),
    .A2(_04050_),
    .A3(_03684_),
    .A4(_03735_),
    .B1(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__a22o_1 _09937_ (.A1(_03692_),
    .A2(_03694_),
    .B1(_03956_),
    .B2(_03959_),
    .X(_04055_));
 sky130_fd_sc_hd__o211ai_1 _09938_ (.A1(_03702_),
    .A2(_03703_),
    .B1(_04019_),
    .C1(_04020_),
    .Y(_04056_));
 sky130_fd_sc_hd__o2111ai_4 _09939_ (.A1(_03635_),
    .A2(_03720_),
    .B1(_01551_),
    .C1(_03730_),
    .D1(_03985_),
    .Y(_04057_));
 sky130_fd_sc_hd__a22o_1 _09940_ (.A1(_00957_),
    .A2(_01540_),
    .B1(_04040_),
    .B2(_04041_),
    .X(_04058_));
 sky130_fd_sc_hd__nand4_1 _09941_ (.A(_01562_),
    .B(_03722_),
    .C(_03730_),
    .D(_04042_),
    .Y(_04060_));
 sky130_fd_sc_hd__o21a_1 _09942_ (.A1(_03732_),
    .A2(_04058_),
    .B1(_04057_),
    .X(_04061_));
 sky130_fd_sc_hd__nand3_1 _09943_ (.A(_04060_),
    .B(_03709_),
    .C(_04057_),
    .Y(_04062_));
 sky130_fd_sc_hd__o211ai_1 _09944_ (.A1(_03732_),
    .A2(_04017_),
    .B1(_04018_),
    .C1(_03710_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand3_1 _09945_ (.A(_04063_),
    .B(_03698_),
    .C(_04062_),
    .Y(_04064_));
 sky130_fd_sc_hd__o211ai_1 _09946_ (.A1(_03710_),
    .A2(_03958_),
    .B1(_03956_),
    .C1(_03699_),
    .Y(_04065_));
 sky130_fd_sc_hd__o221ai_2 _09947_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03710_),
    .B2(_04061_),
    .C1(_04056_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_1 _09948_ (.A(_04055_),
    .B(_04064_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand3_2 _09949_ (.A(_04066_),
    .B(_03687_),
    .C(_04065_),
    .Y(_04068_));
 sky130_fd_sc_hd__o311ai_4 _09950_ (.A1(_03698_),
    .A2(_03789_),
    .A3(_03794_),
    .B1(_03808_),
    .C1(_03882_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand3_1 _09951_ (.A(_04055_),
    .B(_04064_),
    .C(_03672_),
    .Y(_04071_));
 sky130_fd_sc_hd__o221ai_4 _09952_ (.A1(_03666_),
    .A2(_03668_),
    .B1(_03699_),
    .B2(_03807_),
    .C1(_03797_),
    .Y(_04072_));
 sky130_fd_sc_hd__a21oi_1 _09953_ (.A1(_04068_),
    .A2(_04069_),
    .B1(_03653_),
    .Y(_04073_));
 sky130_fd_sc_hd__a21oi_1 _09954_ (.A1(_03643_),
    .A2(_03649_),
    .B1(net32),
    .Y(_04074_));
 sky130_fd_sc_hd__a31oi_4 _09955_ (.A1(_04068_),
    .A2(_04069_),
    .A3(net109),
    .B1(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__o21a_1 _09956_ (.A1(net108),
    .A2(_03733_),
    .B1(net64),
    .X(_04076_));
 sky130_fd_sc_hd__a41oi_4 _09957_ (.A1(_04072_),
    .A2(_03684_),
    .A3(_04071_),
    .A4(_03735_),
    .B1(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__o2bb2ai_1 _09958_ (.A1_N(_04077_),
    .A2_N(_04075_),
    .B1(_04054_),
    .B2(_04051_),
    .Y(_04078_));
 sky130_fd_sc_hd__a211o_1 _09959_ (.A1(net32),
    .A2(_03653_),
    .B1(_04073_),
    .C1(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__o211ai_1 _09960_ (.A1(_04034_),
    .A2(_04031_),
    .B1(_04011_),
    .C1(_04005_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _09961_ (.A(_04036_),
    .B(_04080_),
    .Y(_04082_));
 sky130_fd_sc_hd__a31oi_1 _09962_ (.A1(_04038_),
    .A2(_04078_),
    .A3(_04079_),
    .B1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21oi_1 _09963_ (.A1(_03968_),
    .A2(_03966_),
    .B1(_03952_),
    .Y(_04084_));
 sky130_fd_sc_hd__a22oi_1 _09964_ (.A1(_03965_),
    .A2(_03969_),
    .B1(_04084_),
    .B2(_03950_),
    .Y(_04085_));
 sky130_fd_sc_hd__a211o_1 _09965_ (.A1(_03911_),
    .A2(_03907_),
    .B1(_03929_),
    .C1(_03924_),
    .X(_04086_));
 sky130_fd_sc_hd__o221ai_1 _09966_ (.A1(_03907_),
    .A2(_03911_),
    .B1(_03933_),
    .B2(_04085_),
    .C1(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__o21bai_1 _09967_ (.A1(_03976_),
    .A2(_04083_),
    .B1_N(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__o2bb2ai_1 _09968_ (.A1_N(_04051_),
    .A2_N(_04054_),
    .B1(_04077_),
    .B2(_04075_),
    .Y(_04089_));
 sky130_fd_sc_hd__nor2_1 _09969_ (.A(_04078_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__nand3_1 _09970_ (.A(_03975_),
    .B(_04038_),
    .C(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__o31ai_4 _09971_ (.A1(_03673_),
    .A2(_03681_),
    .A3(_03881_),
    .B1(_03686_),
    .Y(_04093_));
 sky130_fd_sc_hd__o221ai_4 _09972_ (.A1(_03666_),
    .A2(_03668_),
    .B1(_03699_),
    .B2(_03896_),
    .C1(_03899_),
    .Y(_04094_));
 sky130_fd_sc_hd__a2bb2oi_1 _09973_ (.A1_N(_03702_),
    .A2_N(_03703_),
    .B1(_04057_),
    .B2(_04060_),
    .Y(_04095_));
 sky130_fd_sc_hd__o2111a_1 _09974_ (.A1(net114),
    .A2(net110),
    .B1(net62),
    .C1(_05339_),
    .D1(_03734_),
    .X(_04096_));
 sky130_fd_sc_hd__mux4_1 _09975_ (.A0(net63),
    .A1(net62),
    .A2(net31),
    .A3(net30),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04097_));
 sky130_fd_sc_hd__o211a_1 _09976_ (.A1(_03704_),
    .A2(_03706_),
    .B1(net106),
    .C1(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__a31oi_1 _09977_ (.A1(net106),
    .A2(_03957_),
    .A3(_03710_),
    .B1(_03698_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _09978_ (.A(_04021_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__o311ai_2 _09979_ (.A1(_04098_),
    .A2(_03699_),
    .A3(_04095_),
    .B1(_03672_),
    .C1(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand3_2 _09980_ (.A(_04094_),
    .B(_04101_),
    .C(_03658_),
    .Y(_04102_));
 sky130_fd_sc_hd__a21oi_1 _09981_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00088_),
    .Y(_04104_));
 sky130_fd_sc_hd__a31oi_2 _09982_ (.A1(_04102_),
    .A2(net108),
    .A3(_04093_),
    .B1(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__a31o_2 _09983_ (.A1(_04102_),
    .A2(net108),
    .A3(_04093_),
    .B1(_04104_),
    .X(_04106_));
 sky130_fd_sc_hd__a21oi_2 _09984_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00374_),
    .Y(_04107_));
 sky130_fd_sc_hd__a31oi_4 _09985_ (.A1(_04102_),
    .A2(_03735_),
    .A3(_04093_),
    .B1(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__a31o_1 _09986_ (.A1(_04102_),
    .A2(_03735_),
    .A3(_04093_),
    .B1(_04107_),
    .X(_04109_));
 sky130_fd_sc_hd__a31o_1 _09987_ (.A1(_03683_),
    .A2(_03698_),
    .A3(_03835_),
    .B1(_03684_),
    .X(_04110_));
 sky130_fd_sc_hd__o211ai_2 _09988_ (.A1(_03666_),
    .A2(_03668_),
    .B1(_03920_),
    .C1(_03921_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21oi_1 _09989_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03698_),
    .Y(_04112_));
 sky130_fd_sc_hd__o211ai_1 _09990_ (.A1(_03702_),
    .A2(_03703_),
    .B1(net106),
    .C1(_04043_),
    .Y(_04113_));
 sky130_fd_sc_hd__a211o_1 _09991_ (.A1(net30),
    .A2(_03738_),
    .B1(_01562_),
    .C1(_04096_),
    .X(_04115_));
 sky130_fd_sc_hd__o2111a_1 _09992_ (.A1(net114),
    .A2(net110),
    .B1(net61),
    .C1(_05339_),
    .D1(_03734_),
    .X(_04116_));
 sky130_fd_sc_hd__a211o_1 _09993_ (.A1(_03738_),
    .A2(net29),
    .B1(_01551_),
    .C1(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__nand4_1 _09994_ (.A(_04115_),
    .B(_04117_),
    .C(_03709_),
    .D(net106),
    .Y(_04118_));
 sky130_fd_sc_hd__a31o_1 _09995_ (.A1(_04118_),
    .A2(_03698_),
    .A3(_04113_),
    .B1(_03673_),
    .X(_04119_));
 sky130_fd_sc_hd__o211ai_4 _09996_ (.A1(_04112_),
    .A2(_04119_),
    .B1(_03658_),
    .C1(_04111_),
    .Y(_04120_));
 sky130_fd_sc_hd__a21oi_1 _09997_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00385_),
    .Y(_04121_));
 sky130_fd_sc_hd__a31o_1 _09998_ (.A1(_04120_),
    .A2(_03735_),
    .A3(_04110_),
    .B1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__a31oi_2 _09999_ (.A1(_04120_),
    .A2(_03735_),
    .A3(_04110_),
    .B1(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__a21oi_2 _10000_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00099_),
    .Y(_04124_));
 sky130_fd_sc_hd__a31oi_2 _10001_ (.A1(_04120_),
    .A2(net108),
    .A3(_04110_),
    .B1(_04124_),
    .Y(_04126_));
 sky130_fd_sc_hd__a31o_1 _10002_ (.A1(_04120_),
    .A2(net108),
    .A3(_04110_),
    .B1(_04124_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_1 _10003_ (.A(_04123_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a22oi_1 _10004_ (.A1(_04123_),
    .A2(_04127_),
    .B1(_04106_),
    .B2(_04108_),
    .Y(_04129_));
 sky130_fd_sc_hd__o21ai_1 _10005_ (.A1(_04105_),
    .A2(_04109_),
    .B1(_04128_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _10006_ (.A(_04122_),
    .B(_04126_),
    .Y(_04131_));
 sky130_fd_sc_hd__a22oi_1 _10007_ (.A1(_04122_),
    .A2(_04126_),
    .B1(_04109_),
    .B2(_04105_),
    .Y(_04132_));
 sky130_fd_sc_hd__o211ai_1 _10008_ (.A1(_04108_),
    .A2(_04106_),
    .B1(_04131_),
    .C1(_04128_),
    .Y(_04133_));
 sky130_fd_sc_hd__a31o_2 _10009_ (.A1(_03796_),
    .A2(_03698_),
    .A3(_03683_),
    .B1(_03684_),
    .X(_04134_));
 sky130_fd_sc_hd__a21oi_1 _10010_ (.A1(_04062_),
    .A2(_04063_),
    .B1(_03698_),
    .Y(_04135_));
 sky130_fd_sc_hd__a31o_1 _10011_ (.A1(_05339_),
    .A2(_03653_),
    .A3(_03734_),
    .B1(_00066_),
    .X(_04137_));
 sky130_fd_sc_hd__mux4_2 _10012_ (.A0(net61),
    .A1(net60),
    .A2(net29),
    .A3(net28),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04138_));
 sky130_fd_sc_hd__o211ai_2 _10013_ (.A1(_03702_),
    .A2(_03703_),
    .B1(net106),
    .C1(_04097_),
    .Y(_04139_));
 sky130_fd_sc_hd__o211ai_2 _10014_ (.A1(_03704_),
    .A2(_03706_),
    .B1(net106),
    .C1(_04138_),
    .Y(_04140_));
 sky130_fd_sc_hd__a31o_1 _10015_ (.A1(_04139_),
    .A2(_04140_),
    .A3(_03698_),
    .B1(_03673_),
    .X(_04141_));
 sky130_fd_sc_hd__a31oi_2 _10016_ (.A1(_03673_),
    .A2(_03961_),
    .A3(_03962_),
    .B1(_03659_),
    .Y(_04142_));
 sky130_fd_sc_hd__o21ai_2 _10017_ (.A1(_04135_),
    .A2(_04141_),
    .B1(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a21oi_1 _10018_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00066_),
    .Y(_04144_));
 sky130_fd_sc_hd__a31oi_2 _10019_ (.A1(_04143_),
    .A2(net108),
    .A3(_04134_),
    .B1(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a31o_1 _10020_ (.A1(_04143_),
    .A2(net108),
    .A3(_04134_),
    .B1(_04144_),
    .X(_04146_));
 sky130_fd_sc_hd__a21oi_1 _10021_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00352_),
    .Y(_04148_));
 sky130_fd_sc_hd__a31oi_1 _10022_ (.A1(_04143_),
    .A2(_03735_),
    .A3(_04134_),
    .B1(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__a31o_1 _10023_ (.A1(_04143_),
    .A2(_03735_),
    .A3(_04134_),
    .B1(_04148_),
    .X(_04150_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(_04150_),
    .B(_04145_),
    .Y(_04151_));
 sky130_fd_sc_hd__a41o_2 _10025_ (.A1(_03683_),
    .A2(_03698_),
    .A3(_03755_),
    .A4(_03756_),
    .B1(_03684_),
    .X(_04152_));
 sky130_fd_sc_hd__a21oi_1 _10026_ (.A1(_04044_),
    .A2(_04045_),
    .B1(_03698_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand4_1 _10027_ (.A(_03710_),
    .B(_04115_),
    .C(_04117_),
    .D(net106),
    .Y(_04154_));
 sky130_fd_sc_hd__o2111ai_2 _10028_ (.A1(_00352_),
    .A2(_03738_),
    .B1(_04137_),
    .C1(_00957_),
    .D1(_01540_),
    .Y(_04155_));
 sky130_fd_sc_hd__a31o_1 _10029_ (.A1(_05339_),
    .A2(_03653_),
    .A3(_03734_),
    .B1(_00077_),
    .X(_04156_));
 sky130_fd_sc_hd__o221ai_2 _10030_ (.A1(_00946_),
    .A2(_01529_),
    .B1(_03738_),
    .B2(_00363_),
    .C1(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand4_1 _10031_ (.A(_03709_),
    .B(net106),
    .C(_04155_),
    .D(_04157_),
    .Y(_04159_));
 sky130_fd_sc_hd__a31o_1 _10032_ (.A1(_04154_),
    .A2(_04159_),
    .A3(_03698_),
    .B1(_03673_),
    .X(_04160_));
 sky130_fd_sc_hd__a31oi_1 _10033_ (.A1(_03673_),
    .A2(_03944_),
    .A3(_03945_),
    .B1(_03659_),
    .Y(_04161_));
 sky130_fd_sc_hd__o21ai_2 _10034_ (.A1(_04153_),
    .A2(_04160_),
    .B1(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21oi_1 _10035_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00363_),
    .Y(_04163_));
 sky130_fd_sc_hd__a31oi_4 _10036_ (.A1(_04162_),
    .A2(_03735_),
    .A3(_04152_),
    .B1(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__a21oi_1 _10037_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00077_),
    .Y(_04165_));
 sky130_fd_sc_hd__a31o_1 _10038_ (.A1(_04162_),
    .A2(net108),
    .A3(_04152_),
    .B1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__o2bb2ai_1 _10039_ (.A1_N(_04164_),
    .A2_N(_04166_),
    .B1(_04145_),
    .B2(_04150_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand4_1 _10040_ (.A(_04129_),
    .B(_04132_),
    .C(_04151_),
    .D(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o21ai_1 _10041_ (.A1(_04106_),
    .A2(_04108_),
    .B1(_04130_),
    .Y(_04170_));
 sky130_fd_sc_hd__a21oi_1 _10042_ (.A1(_04168_),
    .A2(_04170_),
    .B1(_04091_),
    .Y(_04171_));
 sky130_fd_sc_hd__o21bai_2 _10043_ (.A1(_04171_),
    .A2(_04088_),
    .B1_N(_03878_),
    .Y(_04172_));
 sky130_fd_sc_hd__a31o_2 _10044_ (.A1(_03829_),
    .A2(_03672_),
    .A3(_03682_),
    .B1(_03684_),
    .X(_04173_));
 sky130_fd_sc_hd__mux4_1 _10045_ (.A0(net59),
    .A1(net58),
    .A2(net27),
    .A3(net26),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04174_));
 sky130_fd_sc_hd__nand4_1 _10046_ (.A(_03709_),
    .B(_03722_),
    .C(_03730_),
    .D(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__a311oi_1 _10047_ (.A1(net106),
    .A2(_04138_),
    .A3(_03710_),
    .B1(_03693_),
    .C1(_03691_),
    .Y(_04176_));
 sky130_fd_sc_hd__a21oi_1 _10048_ (.A1(_04176_),
    .A2(_04175_),
    .B1(_03673_),
    .Y(_04177_));
 sky130_fd_sc_hd__o31ai_1 _10049_ (.A1(_03698_),
    .A2(_04095_),
    .A3(_04098_),
    .B1(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a22o_1 _10050_ (.A1(_03667_),
    .A2(_03669_),
    .B1(_04016_),
    .B2(_04024_),
    .X(_04179_));
 sky130_fd_sc_hd__nand3_2 _10051_ (.A(_04179_),
    .B(_03658_),
    .C(_04178_),
    .Y(_04181_));
 sky130_fd_sc_hd__a21oi_1 _10052_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00330_),
    .Y(_04182_));
 sky130_fd_sc_hd__a31oi_2 _10053_ (.A1(_04173_),
    .A2(_04181_),
    .A3(_03735_),
    .B1(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__a31o_2 _10054_ (.A1(_04173_),
    .A2(_04181_),
    .A3(_03735_),
    .B1(_04182_),
    .X(_04184_));
 sky130_fd_sc_hd__a21oi_1 _10055_ (.A1(_03643_),
    .A2(_03649_),
    .B1(_00044_),
    .Y(_04185_));
 sky130_fd_sc_hd__a31oi_2 _10056_ (.A1(_04173_),
    .A2(_04181_),
    .A3(net108),
    .B1(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__a31o_1 _10057_ (.A1(_04173_),
    .A2(_04181_),
    .A3(net108),
    .B1(_04185_),
    .X(_04187_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(_04187_),
    .B(_04183_),
    .Y(_04188_));
 sky130_fd_sc_hd__a21oi_1 _10059_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net55),
    .Y(_04189_));
 sky130_fd_sc_hd__o21ai_1 _10060_ (.A1(net108),
    .A2(_03733_),
    .B1(_00341_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21oi_1 _10061_ (.A1(_03992_),
    .A2(_03994_),
    .B1(_03672_),
    .Y(_04192_));
 sky130_fd_sc_hd__mux4_1 _10062_ (.A0(net58),
    .A1(net55),
    .A2(net26),
    .A3(net23),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04193_));
 sky130_fd_sc_hd__nand3_1 _10063_ (.A(_03699_),
    .B(_04113_),
    .C(_04118_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand4_1 _10064_ (.A(_03709_),
    .B(_03722_),
    .C(_03730_),
    .D(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand4_1 _10065_ (.A(net106),
    .B(_04155_),
    .C(_04157_),
    .D(_03710_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand3_1 _10066_ (.A(_04195_),
    .B(_04196_),
    .C(_03698_),
    .Y(_04197_));
 sky130_fd_sc_hd__a31o_1 _10067_ (.A1(_04194_),
    .A2(_04197_),
    .A3(_03672_),
    .B1(_03659_),
    .X(_04198_));
 sky130_fd_sc_hd__o22a_2 _10068_ (.A1(_03684_),
    .A2(_03844_),
    .B1(_04192_),
    .B2(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__nor2_1 _10069_ (.A(_03736_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__o21ai_1 _10070_ (.A1(_03736_),
    .A2(_04199_),
    .B1(_04190_),
    .Y(_04201_));
 sky130_fd_sc_hd__o21ai_1 _10071_ (.A1(net114),
    .A2(net110),
    .B1(_00055_),
    .Y(_04203_));
 sky130_fd_sc_hd__o21ai_1 _10072_ (.A1(_03653_),
    .A2(_04199_),
    .B1(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21a_2 _10073_ (.A1(_03653_),
    .A2(_04199_),
    .B1(_04203_),
    .X(_04205_));
 sky130_fd_sc_hd__o21ai_1 _10074_ (.A1(_04189_),
    .A2(_04200_),
    .B1(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__a22o_1 _10075_ (.A1(_04187_),
    .A2(_04183_),
    .B1(_04205_),
    .B2(_04201_),
    .X(_04207_));
 sky130_fd_sc_hd__nand2_1 _10076_ (.A(_04184_),
    .B(_04186_),
    .Y(_04208_));
 sky130_fd_sc_hd__o211ai_1 _10077_ (.A1(_03736_),
    .A2(_04199_),
    .B1(_04190_),
    .C1(_04204_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand4_1 _10078_ (.A(_04188_),
    .B(_04206_),
    .C(_04208_),
    .D(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__mux4_1 _10079_ (.A0(net55),
    .A1(net44),
    .A2(net23),
    .A3(net12),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04211_));
 sky130_fd_sc_hd__nand4_1 _10080_ (.A(_03709_),
    .B(_04211_),
    .C(_03730_),
    .D(_03722_),
    .Y(_04212_));
 sky130_fd_sc_hd__a31oi_1 _10081_ (.A1(net106),
    .A2(_04174_),
    .A3(_03710_),
    .B1(_03699_),
    .Y(_04214_));
 sky130_fd_sc_hd__a32oi_2 _10082_ (.A1(_03699_),
    .A2(_04139_),
    .A3(_04140_),
    .B1(_04214_),
    .B2(_04212_),
    .Y(_04215_));
 sky130_fd_sc_hd__or3_1 _10083_ (.A(_03668_),
    .B(_03659_),
    .C(_03666_),
    .X(_04216_));
 sky130_fd_sc_hd__o21a_1 _10084_ (.A1(_04216_),
    .A2(_04215_),
    .B1(_03682_),
    .X(_04217_));
 sky130_fd_sc_hd__o221ai_4 _10085_ (.A1(_04067_),
    .A2(_03672_),
    .B1(_03658_),
    .B2(_03810_),
    .C1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o21ai_1 _10086_ (.A1(net114),
    .A2(net110),
    .B1(net12),
    .Y(_04219_));
 sky130_fd_sc_hd__o21a_2 _10087_ (.A1(_03653_),
    .A2(_04218_),
    .B1(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__inv_2 _10088_ (.A(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a21oi_1 _10089_ (.A1(_03653_),
    .A2(_03734_),
    .B1(net44),
    .Y(_04222_));
 sky130_fd_sc_hd__o311a_2 _10090_ (.A1(_03624_),
    .A2(_03636_),
    .A3(_03638_),
    .B1(_03653_),
    .C1(_04218_),
    .X(_04223_));
 sky130_fd_sc_hd__a21oi_1 _10091_ (.A1(_04218_),
    .A2(_03735_),
    .B1(_04222_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor2_1 _10092_ (.A(_04225_),
    .B(_04220_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21oi_2 _10093_ (.A1(_03653_),
    .A2(_03734_),
    .B1(_00319_),
    .Y(_04227_));
 sky130_fd_sc_hd__a21oi_2 _10094_ (.A1(_04046_),
    .A2(_04047_),
    .B1(_03672_),
    .Y(_04228_));
 sky130_fd_sc_hd__and3_1 _10095_ (.A(_03699_),
    .B(_04154_),
    .C(_04159_),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_1 _10096_ (.A0(net44),
    .A1(net33),
    .A2(net12),
    .A3(net1),
    .S0(_01562_),
    .S1(_03738_),
    .X(_04230_));
 sky130_fd_sc_hd__and3_1 _10097_ (.A(_03709_),
    .B(net106),
    .C(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__a31o_1 _10098_ (.A1(_03710_),
    .A2(_04193_),
    .A3(net106),
    .B1(_03699_),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_1 _10099_ (.A1(_04231_),
    .A2(_04232_),
    .B1(_03672_),
    .Y(_04233_));
 sky130_fd_sc_hd__o21ai_2 _10100_ (.A1(_04229_),
    .A2(_04233_),
    .B1(_03658_),
    .Y(_04234_));
 sky130_fd_sc_hd__a31o_1 _10101_ (.A1(_03783_),
    .A2(_03672_),
    .A3(_03782_),
    .B1(_03658_),
    .X(_04236_));
 sky130_fd_sc_hd__o2111a_1 _10102_ (.A1(_04228_),
    .A2(_04234_),
    .B1(_03735_),
    .C1(_04236_),
    .D1(_03682_),
    .X(_04237_));
 sky130_fd_sc_hd__a21oi_1 _10103_ (.A1(net33),
    .A2(_03736_),
    .B1(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__o2111ai_4 _10104_ (.A1(_04228_),
    .A2(_04234_),
    .B1(net108),
    .C1(_04236_),
    .D1(_03682_),
    .Y(_04239_));
 sky130_fd_sc_hd__o21ai_4 _10105_ (.A1(_00033_),
    .A2(net108),
    .B1(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__o221ai_2 _10106_ (.A1(_00033_),
    .A2(net108),
    .B1(_04227_),
    .B2(_04237_),
    .C1(_04239_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_1 _10107_ (.A(_04220_),
    .B(_04225_),
    .Y(_04242_));
 sky130_fd_sc_hd__a21oi_1 _10108_ (.A1(_04241_),
    .A2(_04242_),
    .B1(_04226_),
    .Y(_04243_));
 sky130_fd_sc_hd__o2bb2ai_1 _10109_ (.A1_N(_04207_),
    .A2_N(_04208_),
    .B1(_04210_),
    .B2(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04164_),
    .B(_04166_),
    .Y(_04245_));
 sky130_fd_sc_hd__a211o_1 _10111_ (.A1(_04145_),
    .A2(_04150_),
    .B1(_04245_),
    .C1(_04167_),
    .X(_04247_));
 sky130_fd_sc_hd__nor2_1 _10112_ (.A(_04091_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a211oi_1 _10113_ (.A1(_04106_),
    .A2(_04108_),
    .B1(_04133_),
    .C1(_03878_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand3_2 _10114_ (.A(_04244_),
    .B(_04248_),
    .C(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand3_1 _10115_ (.A(_03818_),
    .B(_03819_),
    .C(_03870_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21oi_1 _10116_ (.A1(_04251_),
    .A2(_03851_),
    .B1(_03855_),
    .Y(_04252_));
 sky130_fd_sc_hd__o21ai_1 _10117_ (.A1(_03873_),
    .A2(_04252_),
    .B1(_03869_),
    .Y(_04253_));
 sky130_fd_sc_hd__o311a_2 _10118_ (.A1(net109),
    .A2(_03866_),
    .A3(_03862_),
    .B1(_03736_),
    .C1(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__or3b_1 _10119_ (.A(_04227_),
    .B(_04237_),
    .C_N(_04240_),
    .X(_04255_));
 sky130_fd_sc_hd__nand3_4 _10120_ (.A(_04172_),
    .B(_04250_),
    .C(_04254_),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2_1 _10121_ (.A(_03853_),
    .B(net102),
    .Y(_04258_));
 sky130_fd_sc_hd__o21ai_2 _10122_ (.A1(_03759_),
    .A2(net102),
    .B1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(_03834_),
    .A1(_03832_),
    .S(net102),
    .X(_04260_));
 sky130_fd_sc_hd__inv_2 _10124_ (.A(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__mux2_2 _10125_ (.A0(_04030_),
    .A1(_04034_),
    .S(net102),
    .X(_04262_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(_04005_),
    .A1(_04010_),
    .S(net102),
    .X(_04263_));
 sky130_fd_sc_hd__o21ai_1 _10127_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_1 _10128_ (.A(net102),
    .B(_04077_),
    .Y(_04265_));
 sky130_fd_sc_hd__o21ai_2 _10129_ (.A1(_04075_),
    .A2(net102),
    .B1(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2b_1 _10130_ (.A_N(_04054_),
    .B(net101),
    .Y(_04267_));
 sky130_fd_sc_hd__o21ai_1 _10131_ (.A1(_04052_),
    .A2(net101),
    .B1(_04267_),
    .Y(_04269_));
 sky130_fd_sc_hd__or2_1 _10132_ (.A(_03618_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nand2_1 _10133_ (.A(net102),
    .B(_04108_),
    .Y(_04271_));
 sky130_fd_sc_hd__o21ai_1 _10134_ (.A1(_04106_),
    .A2(net101),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__or2_2 _10135_ (.A(_03618_),
    .B(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__nand2_1 _10136_ (.A(_04123_),
    .B(net102),
    .Y(_04274_));
 sky130_fd_sc_hd__o21a_1 _10137_ (.A1(_04127_),
    .A2(net101),
    .B1(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__o221a_1 _10138_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04127_),
    .B2(net101),
    .C1(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__nand2_1 _10139_ (.A(net101),
    .B(_04238_),
    .Y(_04277_));
 sky130_fd_sc_hd__a31o_1 _10140_ (.A1(_04172_),
    .A2(_04250_),
    .A3(_04254_),
    .B1(_04238_),
    .X(_04278_));
 sky130_fd_sc_hd__nand4_2 _10141_ (.A(_04172_),
    .B(_04240_),
    .C(_04250_),
    .D(_04254_),
    .Y(_04280_));
 sky130_fd_sc_hd__o22a_1 _10142_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04240_),
    .B2(net101),
    .X(_04281_));
 sky130_fd_sc_hd__o211ai_4 _10143_ (.A1(_04240_),
    .A2(net101),
    .B1(_03617_),
    .C1(_04277_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_1 _10144_ (.A(_04225_),
    .B(net101),
    .Y(_04283_));
 sky130_fd_sc_hd__o21ai_2 _10145_ (.A1(_04222_),
    .A2(_04223_),
    .B1(net101),
    .Y(_04284_));
 sky130_fd_sc_hd__o21ai_1 _10146_ (.A1(_04221_),
    .A2(net101),
    .B1(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__o21ai_1 _10147_ (.A1(_04220_),
    .A2(net101),
    .B1(_04283_),
    .Y(_04286_));
 sky130_fd_sc_hd__nand2_1 _10148_ (.A(_04282_),
    .B(_04285_),
    .Y(_04287_));
 sky130_fd_sc_hd__o221ai_4 _10149_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04221_),
    .B2(net101),
    .C1(_04284_),
    .Y(_04288_));
 sky130_fd_sc_hd__o2111ai_4 _10150_ (.A1(_04256_),
    .A2(_04220_),
    .B1(_04280_),
    .C1(_04278_),
    .D1(_04283_),
    .Y(_04289_));
 sky130_fd_sc_hd__o21ai_2 _10151_ (.A1(_04189_),
    .A2(_04200_),
    .B1(net101),
    .Y(_04291_));
 sky130_fd_sc_hd__o21ai_2 _10152_ (.A1(_04205_),
    .A2(net101),
    .B1(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__o211ai_4 _10153_ (.A1(_04205_),
    .A2(net101),
    .B1(_03617_),
    .C1(_04291_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand3_2 _10154_ (.A(_04282_),
    .B(_04288_),
    .C(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(net101),
    .B(_04183_),
    .Y(_04295_));
 sky130_fd_sc_hd__o21ai_2 _10156_ (.A1(_04187_),
    .A2(net101),
    .B1(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21a_1 _10157_ (.A1(_04187_),
    .A2(net101),
    .B1(_04295_),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_04164_),
    .B(net101),
    .Y(_04298_));
 sky130_fd_sc_hd__o21ai_1 _10159_ (.A1(_04166_),
    .A2(net101),
    .B1(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__o21a_1 _10160_ (.A1(_04166_),
    .A2(net101),
    .B1(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_1 _10161_ (.A(net101),
    .B(_04149_),
    .Y(_04302_));
 sky130_fd_sc_hd__o21ai_2 _10162_ (.A1(_04146_),
    .A2(net101),
    .B1(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__o21a_1 _10163_ (.A1(_04146_),
    .A2(net101),
    .B1(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__nand3_2 _10164_ (.A(_04296_),
    .B(_04299_),
    .C(_04303_),
    .Y(_04305_));
 sky130_fd_sc_hd__o21ai_1 _10165_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04300_),
    .Y(_04306_));
 sky130_fd_sc_hd__o221a_1 _10166_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04187_),
    .B2(net101),
    .C1(_04295_),
    .X(_04307_));
 sky130_fd_sc_hd__a21oi_1 _10167_ (.A1(_04305_),
    .A2(_03617_),
    .B1(_04294_),
    .Y(_04308_));
 sky130_fd_sc_hd__a211oi_4 _10168_ (.A1(_04305_),
    .A2(_03617_),
    .B1(_04276_),
    .C1(_04294_),
    .Y(_04309_));
 sky130_fd_sc_hd__o2111a_1 _10169_ (.A1(_04266_),
    .A2(_03618_),
    .B1(_04273_),
    .C1(_04270_),
    .D1(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__o2111ai_2 _10170_ (.A1(_04266_),
    .A2(_03618_),
    .B1(_04273_),
    .C1(_04270_),
    .D1(_04309_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21o_1 _10171_ (.A1(_03617_),
    .A2(_04263_),
    .B1(_04311_),
    .X(_04313_));
 sky130_fd_sc_hd__o211ai_1 _10172_ (.A1(_03618_),
    .A2(_04262_),
    .B1(_04264_),
    .C1(_04310_),
    .Y(_04314_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(_03952_),
    .A1(_03950_),
    .S(net102),
    .X(_04315_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(_03968_),
    .A1(_03965_),
    .S(net102),
    .X(_04316_));
 sky130_fd_sc_hd__a41o_1 _10175_ (.A1(_04262_),
    .A2(_04310_),
    .A3(_04315_),
    .A4(_04264_),
    .B1(_03618_),
    .X(_04317_));
 sky130_fd_sc_hd__o21ai_1 _10176_ (.A1(_03618_),
    .A2(_04316_),
    .B1(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(_03924_),
    .A1(_03928_),
    .S(net102),
    .X(_04319_));
 sky130_fd_sc_hd__o211ai_2 _10178_ (.A1(_03618_),
    .A2(_04316_),
    .B1(_04319_),
    .C1(_04317_),
    .Y(_04320_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(_03908_),
    .A1(_03911_),
    .S(net102),
    .X(_04321_));
 sky130_fd_sc_hd__o21ai_1 _10180_ (.A1(_04320_),
    .A2(_04321_),
    .B1(_03617_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _10181_ (.A(_03788_),
    .B(net102),
    .Y(_04324_));
 sky130_fd_sc_hd__o21ai_1 _10182_ (.A1(_03786_),
    .A2(net102),
    .B1(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(_03814_),
    .A1(_03812_),
    .S(net102),
    .X(_04326_));
 sky130_fd_sc_hd__o21ai_2 _10184_ (.A1(_03618_),
    .A2(_04325_),
    .B1(_04322_),
    .Y(_04327_));
 sky130_fd_sc_hd__a21oi_1 _10185_ (.A1(_03617_),
    .A2(_04326_),
    .B1(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(_03846_),
    .A1(_03848_),
    .S(net102),
    .X(_04329_));
 sky130_fd_sc_hd__o31a_2 _10187_ (.A1(_04326_),
    .A2(_04329_),
    .A3(_04327_),
    .B1(_03617_),
    .X(_04330_));
 sky130_fd_sc_hd__a21oi_1 _10188_ (.A1(_03617_),
    .A2(_04261_),
    .B1(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_1 _10189_ (.A(net102),
    .B(_03857_),
    .Y(_04332_));
 sky130_fd_sc_hd__o21a_1 _10190_ (.A1(_03859_),
    .A2(net102),
    .B1(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__o31a_1 _10191_ (.A1(_04259_),
    .A2(_04261_),
    .A3(_04330_),
    .B1(_03617_),
    .X(_04335_));
 sky130_fd_sc_hd__o41a_1 _10192_ (.A1(_04259_),
    .A2(_04261_),
    .A3(_04333_),
    .A4(_04330_),
    .B1(_03617_),
    .X(_04336_));
 sky130_fd_sc_hd__mux2_1 _10193_ (.A0(_03863_),
    .A1(_03866_),
    .S(net102),
    .X(_04337_));
 sky130_fd_sc_hd__a211o_1 _10194_ (.A1(_04333_),
    .A2(_03617_),
    .B1(_04337_),
    .C1(_04335_),
    .X(_04338_));
 sky130_fd_sc_hd__a311oi_1 _10195_ (.A1(_00000_),
    .A2(_00836_),
    .A3(_00847_),
    .B1(net109),
    .C1(net102),
    .Y(_04339_));
 sky130_fd_sc_hd__a31o_1 _10196_ (.A1(_00792_),
    .A2(_03736_),
    .A3(net102),
    .B1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__o311a_1 _10197_ (.A1(_04337_),
    .A2(_04333_),
    .A3(_04335_),
    .B1(_04340_),
    .C1(_03617_),
    .X(_04341_));
 sky130_fd_sc_hd__a21oi_2 _10198_ (.A1(_04338_),
    .A2(_03617_),
    .B1(_04340_),
    .Y(_04342_));
 sky130_fd_sc_hd__nor2_1 _10199_ (.A(_04341_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__or3b_1 _10200_ (.A(_00869_),
    .B(net109),
    .C_N(net102),
    .X(_04344_));
 sky130_fd_sc_hd__o31a_1 _10201_ (.A1(_00781_),
    .A2(_03735_),
    .A3(net102),
    .B1(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__or3_2 _10202_ (.A(_04341_),
    .B(_04342_),
    .C(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _10203_ (.A(_04336_),
    .B(_04337_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_04338_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _10205_ (.A(_03863_),
    .B(net102),
    .Y(_04350_));
 sky130_fd_sc_hd__o31a_2 _10206_ (.A1(_03864_),
    .A2(_03865_),
    .A3(net102),
    .B1(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__nor2_1 _10207_ (.A(_04349_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__o311a_1 _10208_ (.A1(_04259_),
    .A2(_04261_),
    .A3(_04330_),
    .B1(_04333_),
    .C1(_03617_),
    .X(_04353_));
 sky130_fd_sc_hd__nor2_1 _10209_ (.A(_04333_),
    .B(_04335_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_03859_),
    .B(net102),
    .Y(_04355_));
 sky130_fd_sc_hd__o21a_1 _10211_ (.A1(_03857_),
    .A2(net102),
    .B1(_04355_),
    .X(_04357_));
 sky130_fd_sc_hd__nor3_1 _10212_ (.A(_04353_),
    .B(_04354_),
    .C(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__xor2_1 _10213_ (.A(_04259_),
    .B(_04331_),
    .X(_04359_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(_03853_),
    .B(net102),
    .Y(_04360_));
 sky130_fd_sc_hd__a21o_1 _10215_ (.A1(_03759_),
    .A2(net102),
    .B1(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__nor2_1 _10216_ (.A(_04359_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__a211o_1 _10217_ (.A1(_03759_),
    .A2(net102),
    .B1(_04360_),
    .C1(_04359_),
    .X(_04363_));
 sky130_fd_sc_hd__xor2_1 _10218_ (.A(_04260_),
    .B(_04330_),
    .X(_04364_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(_03832_),
    .A1(_03834_),
    .S(net102),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _10220_ (.A(_04364_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__xor2_1 _10221_ (.A(_04328_),
    .B(_04329_),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(_03848_),
    .A1(_03846_),
    .S(net102),
    .X(_04369_));
 sky130_fd_sc_hd__and2b_1 _10223_ (.A_N(_04368_),
    .B(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(_03812_),
    .A1(_03814_),
    .S(net102),
    .X(_04371_));
 sky130_fd_sc_hd__xor2_1 _10225_ (.A(_04326_),
    .B(_04327_),
    .X(_04372_));
 sky130_fd_sc_hd__and2_1 _10226_ (.A(_04372_),
    .B(_04371_),
    .X(_04373_));
 sky130_fd_sc_hd__nor2_1 _10227_ (.A(_04371_),
    .B(_04372_),
    .Y(_04374_));
 sky130_fd_sc_hd__or2_2 _10228_ (.A(_04373_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__inv_2 _10229_ (.A(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__xnor2_1 _10230_ (.A(_04322_),
    .B(_04325_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _10231_ (.A(_03786_),
    .B(net102),
    .Y(_04379_));
 sky130_fd_sc_hd__o21ai_1 _10232_ (.A1(_03788_),
    .A2(net102),
    .B1(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__and2b_1 _10233_ (.A_N(_04377_),
    .B(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__and3_1 _10234_ (.A(_04320_),
    .B(_04321_),
    .C(_03617_),
    .X(_04382_));
 sky130_fd_sc_hd__a21oi_1 _10235_ (.A1(_04320_),
    .A2(_03617_),
    .B1(_04321_),
    .Y(_04383_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(_03911_),
    .A1(_03908_),
    .S(net102),
    .X(_04384_));
 sky130_fd_sc_hd__inv_2 _10237_ (.A(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__nor3_1 _10238_ (.A(_04382_),
    .B(_04383_),
    .C(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__xor2_1 _10239_ (.A(_04318_),
    .B(_04319_),
    .X(_04387_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(_03928_),
    .A1(_03924_),
    .S(net102),
    .X(_04388_));
 sky130_fd_sc_hd__nor2_1 _10241_ (.A(_04388_),
    .B(_04387_),
    .Y(_04390_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(_03965_),
    .A1(_03968_),
    .S(net102),
    .X(_04391_));
 sky130_fd_sc_hd__xnor2_1 _10243_ (.A(_04316_),
    .B(_04317_),
    .Y(_04392_));
 sky130_fd_sc_hd__nor2_1 _10244_ (.A(_04391_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__and2_1 _10245_ (.A(_04392_),
    .B(_04391_),
    .X(_04394_));
 sky130_fd_sc_hd__nor2_2 _10246_ (.A(_04393_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__xor2_1 _10247_ (.A(_04314_),
    .B(_04315_),
    .X(_04396_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(_03950_),
    .A1(_03952_),
    .S(net102),
    .X(_04397_));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__or2_1 _10250_ (.A(_04397_),
    .B(_04396_),
    .X(_04399_));
 sky130_fd_sc_hd__xor2_4 _10251_ (.A(_04262_),
    .B(_04313_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_2 _10252_ (.A0(_04034_),
    .A1(_04030_),
    .S(net102),
    .X(_04402_));
 sky130_fd_sc_hd__xor2_2 _10253_ (.A(_04401_),
    .B(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__nor2_1 _10254_ (.A(_04263_),
    .B(_04311_),
    .Y(_04404_));
 sky130_fd_sc_hd__and2_1 _10255_ (.A(_04263_),
    .B(_04311_),
    .X(_04405_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(_04010_),
    .A1(_04005_),
    .S(net102),
    .X(_04406_));
 sky130_fd_sc_hd__o21bai_1 _10257_ (.A1(_04404_),
    .A2(_04405_),
    .B1_N(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__or3b_1 _10258_ (.A(_04404_),
    .B(_04405_),
    .C_N(_04406_),
    .X(_04408_));
 sky130_fd_sc_hd__and4_1 _10259_ (.A(_04270_),
    .B(_04309_),
    .C(_04273_),
    .D(_04266_),
    .X(_04409_));
 sky130_fd_sc_hd__a31oi_1 _10260_ (.A1(_04309_),
    .A2(_04273_),
    .A3(_04270_),
    .B1(_04266_),
    .Y(_04410_));
 sky130_fd_sc_hd__or2_1 _10261_ (.A(_04409_),
    .B(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__nand2_1 _10262_ (.A(_04075_),
    .B(net102),
    .Y(_04413_));
 sky130_fd_sc_hd__o21a_1 _10263_ (.A1(_04077_),
    .A2(net102),
    .B1(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__o221a_1 _10264_ (.A1(net102),
    .A2(_04077_),
    .B1(_04410_),
    .B2(_04409_),
    .C1(_04413_),
    .X(_04415_));
 sky130_fd_sc_hd__inv_2 _10265_ (.A(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor2_1 _10266_ (.A(_04414_),
    .B(_04412_),
    .Y(_04417_));
 sky130_fd_sc_hd__o2111a_1 _10267_ (.A1(_04052_),
    .A2(net101),
    .B1(_04267_),
    .C1(_04273_),
    .D1(_04309_),
    .X(_04418_));
 sky130_fd_sc_hd__a21boi_1 _10268_ (.A1(_04309_),
    .A2(_04273_),
    .B1_N(_04269_),
    .Y(_04419_));
 sky130_fd_sc_hd__or2_1 _10269_ (.A(_04418_),
    .B(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _10270_ (.A(_04418_),
    .B(_04419_),
    .Y(_04421_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(_04054_),
    .A1(_04052_),
    .S(net101),
    .X(_04423_));
 sky130_fd_sc_hd__inv_2 _10272_ (.A(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__or3_1 _10273_ (.A(_04418_),
    .B(_04423_),
    .C(_04419_),
    .X(_04425_));
 sky130_fd_sc_hd__o21ai_1 _10274_ (.A1(_04418_),
    .A2(_04419_),
    .B1(_04423_),
    .Y(_04426_));
 sky130_fd_sc_hd__o211a_1 _10275_ (.A1(_04106_),
    .A2(net101),
    .B1(_04271_),
    .C1(_04309_),
    .X(_04427_));
 sky130_fd_sc_hd__and2b_1 _10276_ (.A_N(_04309_),
    .B(_04272_),
    .X(_04428_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(_04108_),
    .A1(_04105_),
    .S(net102),
    .X(_04429_));
 sky130_fd_sc_hd__or3b_1 _10278_ (.A(_04427_),
    .B(_04428_),
    .C_N(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__o21bai_1 _10279_ (.A1(_04427_),
    .A2(_04428_),
    .B1_N(_04429_),
    .Y(_04431_));
 sky130_fd_sc_hd__nor2_1 _10280_ (.A(_04275_),
    .B(_04308_),
    .Y(_04432_));
 sky130_fd_sc_hd__o211a_1 _10281_ (.A1(_04127_),
    .A2(net101),
    .B1(_04274_),
    .C1(_04308_),
    .X(_04434_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_04308_),
    .B(_04275_),
    .Y(_04435_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(_04123_),
    .A1(_04126_),
    .S(net102),
    .X(_04436_));
 sky130_fd_sc_hd__o21bai_1 _10284_ (.A1(_04432_),
    .A2(_04434_),
    .B1_N(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand4_4 _10285_ (.A(_04282_),
    .B(_04288_),
    .C(_04293_),
    .D(_04296_),
    .Y(_04438_));
 sky130_fd_sc_hd__a21oi_1 _10286_ (.A1(_04289_),
    .A2(_03617_),
    .B1(_04307_),
    .Y(_04439_));
 sky130_fd_sc_hd__o211ai_1 _10287_ (.A1(_04300_),
    .A2(_04438_),
    .B1(_04304_),
    .C1(_03617_),
    .Y(_04440_));
 sky130_fd_sc_hd__o2111ai_1 _10288_ (.A1(_03618_),
    .A2(_04292_),
    .B1(_04303_),
    .C1(_04306_),
    .D1(_04439_),
    .Y(_04441_));
 sky130_fd_sc_hd__o211ai_1 _10289_ (.A1(_04300_),
    .A2(_04438_),
    .B1(_04303_),
    .C1(_03617_),
    .Y(_04442_));
 sky130_fd_sc_hd__nand4_1 _10290_ (.A(_04439_),
    .B(_04306_),
    .C(_04304_),
    .D(_04293_),
    .Y(_04443_));
 sky130_fd_sc_hd__mux2_1 _10291_ (.A0(_04150_),
    .A1(_04146_),
    .S(net101),
    .X(_04445_));
 sky130_fd_sc_hd__inv_2 _10292_ (.A(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand3_1 _10293_ (.A(_04440_),
    .B(_04441_),
    .C(_04445_),
    .Y(_04447_));
 sky130_fd_sc_hd__inv_2 _10294_ (.A(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand3_1 _10295_ (.A(_04442_),
    .B(_04443_),
    .C(_04446_),
    .Y(_04449_));
 sky130_fd_sc_hd__and2_1 _10296_ (.A(_04447_),
    .B(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__a21o_1 _10297_ (.A1(_04439_),
    .A2(_04293_),
    .B1(_04299_),
    .X(_04451_));
 sky130_fd_sc_hd__a21o_1 _10298_ (.A1(_04438_),
    .A2(_03617_),
    .B1(_04300_),
    .X(_04452_));
 sky130_fd_sc_hd__nand2_1 _10299_ (.A(_04166_),
    .B(net101),
    .Y(_04453_));
 sky130_fd_sc_hd__o21ai_1 _10300_ (.A1(_04164_),
    .A2(net101),
    .B1(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21o_2 _10301_ (.A1(_04451_),
    .A2(_04452_),
    .B1(_04454_),
    .X(_04456_));
 sky130_fd_sc_hd__nand3_2 _10302_ (.A(_04451_),
    .B(_04452_),
    .C(_04454_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2_2 _10303_ (.A(_04294_),
    .B(_04297_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand2_1 _10304_ (.A(_04438_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__nor2_1 _10305_ (.A(_04184_),
    .B(net101),
    .Y(_04460_));
 sky130_fd_sc_hd__and2_1 _10306_ (.A(net101),
    .B(_04186_),
    .X(_04461_));
 sky130_fd_sc_hd__nand2_1 _10307_ (.A(net101),
    .B(_04186_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21ai_2 _10308_ (.A1(_04184_),
    .A2(net101),
    .B1(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__o2111ai_4 _10309_ (.A1(_04184_),
    .A2(net101),
    .B1(_04438_),
    .C1(_04458_),
    .D1(_04462_),
    .Y(_04464_));
 sky130_fd_sc_hd__o2bb2ai_2 _10310_ (.A1_N(_04438_),
    .A2_N(_04458_),
    .B1(_04460_),
    .B2(_04461_),
    .Y(_04465_));
 sky130_fd_sc_hd__nand3b_1 _10311_ (.A_N(_04292_),
    .B(_03617_),
    .C(_04289_),
    .Y(_04467_));
 sky130_fd_sc_hd__o211ai_1 _10312_ (.A1(_03618_),
    .A2(_04285_),
    .B1(_04292_),
    .C1(_04282_),
    .Y(_04468_));
 sky130_fd_sc_hd__a21o_1 _10313_ (.A1(_04289_),
    .A2(_03617_),
    .B1(_04292_),
    .X(_04469_));
 sky130_fd_sc_hd__o211ai_1 _10314_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_04292_),
    .C1(_04289_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _10315_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__o21ai_1 _10316_ (.A1(net23),
    .A2(net108),
    .B1(net101),
    .Y(_04472_));
 sky130_fd_sc_hd__o21ai_2 _10317_ (.A1(_04201_),
    .A2(net101),
    .B1(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21o_1 _10318_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__nand3_1 _10319_ (.A(_04467_),
    .B(_04468_),
    .C(_04473_),
    .Y(_04475_));
 sky130_fd_sc_hd__o2111ai_1 _10320_ (.A1(_04240_),
    .A2(net101),
    .B1(_03617_),
    .C1(_04277_),
    .D1(_04286_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21oi_1 _10321_ (.A1(_04281_),
    .A2(_04277_),
    .B1(_04285_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand2_1 _10322_ (.A(_04287_),
    .B(_04476_),
    .Y(_04479_));
 sky130_fd_sc_hd__o311a_1 _10323_ (.A1(net110),
    .A2(net114),
    .A3(_04218_),
    .B1(_04219_),
    .C1(net101),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_1 _10324_ (.A(_04225_),
    .B(net101),
    .Y(_04481_));
 sky130_fd_sc_hd__a21o_1 _10325_ (.A1(_04220_),
    .A2(net101),
    .B1(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__o22ai_2 _10326_ (.A1(_04480_),
    .A2(_04481_),
    .B1(_04282_),
    .B2(_04286_),
    .Y(_04483_));
 sky130_fd_sc_hd__nor2_1 _10327_ (.A(_04482_),
    .B(_04479_),
    .Y(_04484_));
 sky130_fd_sc_hd__o21a_1 _10328_ (.A1(_04227_),
    .A2(_04237_),
    .B1(_04240_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _10329_ (.A(_04241_),
    .B(_04255_),
    .Y(_04486_));
 sky130_fd_sc_hd__and2_1 _10330_ (.A(_04486_),
    .B(net65),
    .X(_04487_));
 sky130_fd_sc_hd__a21oi_1 _10331_ (.A1(_04486_),
    .A2(net65),
    .B1(_04485_),
    .Y(_04489_));
 sky130_fd_sc_hd__o22ai_2 _10332_ (.A1(_04485_),
    .A2(_04487_),
    .B1(_04478_),
    .B2(_04483_),
    .Y(_04490_));
 sky130_fd_sc_hd__o31a_1 _10333_ (.A1(_04480_),
    .A2(_04481_),
    .A3(_04479_),
    .B1(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__o211ai_2 _10334_ (.A1(_04482_),
    .A2(_04479_),
    .B1(_04475_),
    .C1(_04490_),
    .Y(_04492_));
 sky130_fd_sc_hd__o2111ai_4 _10335_ (.A1(_04473_),
    .A2(_04471_),
    .B1(_04465_),
    .C1(_04464_),
    .D1(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__o31a_1 _10336_ (.A1(_04459_),
    .A2(_04460_),
    .A3(_04461_),
    .B1(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__o211ai_4 _10337_ (.A1(_04463_),
    .A2(_04459_),
    .B1(_04457_),
    .C1(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__and3_1 _10338_ (.A(_04495_),
    .B(_04450_),
    .C(_04456_),
    .X(_04496_));
 sky130_fd_sc_hd__a31oi_4 _10339_ (.A1(_04495_),
    .A2(_04450_),
    .A3(_04456_),
    .B1(_04448_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand3b_1 _10340_ (.A_N(_04432_),
    .B(_04435_),
    .C(_04436_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _10341_ (.A(_04437_),
    .B(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__o21ai_1 _10342_ (.A1(_04500_),
    .A2(_04497_),
    .B1(_04437_),
    .Y(_04501_));
 sky130_fd_sc_hd__o211ai_1 _10343_ (.A1(_04500_),
    .A2(_04497_),
    .B1(_04437_),
    .C1(_04431_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _10344_ (.A(_04430_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__o2bb2ai_1 _10345_ (.A1_N(_04430_),
    .A2_N(_04502_),
    .B1(_04421_),
    .B2(_04424_),
    .Y(_04504_));
 sky130_fd_sc_hd__o21ai_1 _10346_ (.A1(_04420_),
    .A2(_04423_),
    .B1(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__o211ai_1 _10347_ (.A1(_04423_),
    .A2(_04420_),
    .B1(_04416_),
    .C1(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__a31o_1 _10348_ (.A1(_04416_),
    .A2(_04425_),
    .A3(_04504_),
    .B1(_04417_),
    .X(_04507_));
 sky130_fd_sc_hd__o211ai_1 _10349_ (.A1(_04414_),
    .A2(_04412_),
    .B1(_04408_),
    .C1(_04506_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_1 _10350_ (.A(_04407_),
    .B(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand3_1 _10351_ (.A(_04508_),
    .B(_04403_),
    .C(_04407_),
    .Y(_04511_));
 sky130_fd_sc_hd__o21ai_2 _10352_ (.A1(_04401_),
    .A2(_04402_),
    .B1(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__o211ai_2 _10353_ (.A1(_04402_),
    .A2(_04401_),
    .B1(_04399_),
    .C1(_04511_),
    .Y(_04513_));
 sky130_fd_sc_hd__a21bo_1 _10354_ (.A1(_04398_),
    .A2(_04512_),
    .B1_N(_04399_),
    .X(_04514_));
 sky130_fd_sc_hd__a31oi_2 _10355_ (.A1(_04513_),
    .A2(_04395_),
    .A3(_04398_),
    .B1(_04393_),
    .Y(_04515_));
 sky130_fd_sc_hd__a31o_1 _10356_ (.A1(_04513_),
    .A2(_04395_),
    .A3(_04398_),
    .B1(_04393_),
    .X(_04516_));
 sky130_fd_sc_hd__nand2_1 _10357_ (.A(_04387_),
    .B(_04388_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand2b_1 _10358_ (.A_N(_04390_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_1 _10359_ (.A1(_04516_),
    .A2(_04517_),
    .B1(_04390_),
    .Y(_04519_));
 sky130_fd_sc_hd__o21bai_2 _10360_ (.A1(_04518_),
    .A2(_04515_),
    .B1_N(_04390_),
    .Y(_04520_));
 sky130_fd_sc_hd__o21a_1 _10361_ (.A1(_04382_),
    .A2(_04383_),
    .B1(_04385_),
    .X(_04522_));
 sky130_fd_sc_hd__or2_1 _10362_ (.A(_04386_),
    .B(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__inv_2 _10363_ (.A(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__a21oi_2 _10364_ (.A1(_04520_),
    .A2(_04524_),
    .B1(_04386_),
    .Y(_04525_));
 sky130_fd_sc_hd__o32ai_1 _10365_ (.A1(_04382_),
    .A2(_04383_),
    .A3(_04385_),
    .B1(_04523_),
    .B2(_04519_),
    .Y(_04526_));
 sky130_fd_sc_hd__and2b_1 _10366_ (.A_N(_04380_),
    .B(_04377_),
    .X(_04527_));
 sky130_fd_sc_hd__or2_2 _10367_ (.A(_04381_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__inv_2 _10368_ (.A(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__a21oi_1 _10369_ (.A1(_04526_),
    .A2(_04529_),
    .B1(_04381_),
    .Y(_04530_));
 sky130_fd_sc_hd__o21bai_2 _10370_ (.A1(_04528_),
    .A2(_04525_),
    .B1_N(_04381_),
    .Y(_04531_));
 sky130_fd_sc_hd__a21oi_1 _10371_ (.A1(_04531_),
    .A2(_04376_),
    .B1(_04373_),
    .Y(_04533_));
 sky130_fd_sc_hd__o21bai_1 _10372_ (.A1(_04375_),
    .A2(_04530_),
    .B1_N(_04373_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2b_1 _10373_ (.A_N(_04369_),
    .B(_04368_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2b_1 _10374_ (.A_N(_04370_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__a21oi_1 _10375_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04370_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21bai_2 _10376_ (.A1(_04536_),
    .A2(_04533_),
    .B1_N(_04370_),
    .Y(_04538_));
 sky130_fd_sc_hd__and2_1 _10377_ (.A(_04364_),
    .B(_04365_),
    .X(_04539_));
 sky130_fd_sc_hd__or2_1 _10378_ (.A(_04366_),
    .B(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__inv_2 _10379_ (.A(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21oi_2 _10380_ (.A1(_04538_),
    .A2(_04541_),
    .B1(_04366_),
    .Y(_04542_));
 sky130_fd_sc_hd__o21bai_1 _10381_ (.A1(_04540_),
    .A2(_04537_),
    .B1_N(_04366_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_04359_),
    .B(_04361_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_2 _10383_ (.A(_04363_),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__inv_2 _10384_ (.A(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand2_1 _10385_ (.A(_04544_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__a21oi_1 _10386_ (.A1(_04544_),
    .A2(_04547_),
    .B1(_04362_),
    .Y(_04549_));
 sky130_fd_sc_hd__o21bai_1 _10387_ (.A1(_04546_),
    .A2(_04542_),
    .B1_N(_04362_),
    .Y(_04550_));
 sky130_fd_sc_hd__o21a_1 _10388_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04357_),
    .X(_04551_));
 sky130_fd_sc_hd__or2_2 _10389_ (.A(_04358_),
    .B(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__inv_2 _10390_ (.A(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21oi_1 _10391_ (.A1(_04363_),
    .A2(_04548_),
    .B1(_04552_),
    .Y(_04555_));
 sky130_fd_sc_hd__a21oi_1 _10392_ (.A1(_04550_),
    .A2(_04553_),
    .B1(_04358_),
    .Y(_04556_));
 sky130_fd_sc_hd__o32ai_2 _10393_ (.A1(_04353_),
    .A2(_04354_),
    .A3(_04357_),
    .B1(_04552_),
    .B2(_04549_),
    .Y(_04557_));
 sky130_fd_sc_hd__and2_1 _10394_ (.A(_04349_),
    .B(_04351_),
    .X(_04558_));
 sky130_fd_sc_hd__or2_1 _10395_ (.A(_04352_),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__inv_2 _10396_ (.A(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_2 _10397_ (.A(_04557_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__a21oi_1 _10398_ (.A1(_04557_),
    .A2(_04560_),
    .B1(_04352_),
    .Y(_04562_));
 sky130_fd_sc_hd__o21bai_1 _10399_ (.A1(_04559_),
    .A2(_04556_),
    .B1_N(_04352_),
    .Y(_04563_));
 sky130_fd_sc_hd__o311a_1 _10400_ (.A1(_00781_),
    .A2(net102),
    .A3(_03735_),
    .B1(_04344_),
    .C1(_04343_),
    .X(_04564_));
 sky130_fd_sc_hd__nor2_1 _10401_ (.A(_04346_),
    .B(_04343_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_2 _10402_ (.A(_04564_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o21ai_4 _10403_ (.A1(_04564_),
    .A2(_04566_),
    .B1(_04563_),
    .Y(_04568_));
 sky130_fd_sc_hd__o32ai_4 _10404_ (.A1(_04341_),
    .A2(_04342_),
    .A3(_04346_),
    .B1(_04567_),
    .B2(_04562_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_2 _10405_ (.A(_04338_),
    .B(_04340_),
    .Y(_04570_));
 sky130_fd_sc_hd__inv_2 _10406_ (.A(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__a22oi_4 _10407_ (.A1(_03617_),
    .A2(_04571_),
    .B1(_04568_),
    .B2(_04347_),
    .Y(_04572_));
 sky130_fd_sc_hd__o21ai_4 _10408_ (.A1(_03618_),
    .A2(_04570_),
    .B1(_04569_),
    .Y(_04573_));
 sky130_fd_sc_hd__o21bai_1 _10409_ (.A1(_04478_),
    .A2(_04483_),
    .B1_N(_04484_),
    .Y(_04574_));
 sky130_fd_sc_hd__xor2_2 _10410_ (.A(_04489_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__inv_2 _10411_ (.A(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__a221o_1 _10412_ (.A1(_03617_),
    .A2(_04571_),
    .B1(_04568_),
    .B2(_04347_),
    .C1(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__nor2_1 _10413_ (.A(net65),
    .B(_04486_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor2_1 _10414_ (.A(_04487_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__inv_2 _10415_ (.A(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o211ai_4 _10416_ (.A1(_04349_),
    .A2(_04351_),
    .B1(_04561_),
    .C1(_04567_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_8 _10417_ (.A(_04568_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__o31ai_1 _10418_ (.A1(_04581_),
    .A2(_04583_),
    .A3(_04572_),
    .B1(_04578_),
    .Y(_04584_));
 sky130_fd_sc_hd__xnor2_2 _10419_ (.A(_04542_),
    .B(_04546_),
    .Y(_04585_));
 sky130_fd_sc_hd__a211o_1 _10420_ (.A1(_04550_),
    .A2(_04553_),
    .B1(_04560_),
    .C1(_04358_),
    .X(_04586_));
 sky130_fd_sc_hd__and3_1 _10421_ (.A(_04363_),
    .B(_04548_),
    .C(_04552_),
    .X(_04588_));
 sky130_fd_sc_hd__nor2_2 _10422_ (.A(_04555_),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__xnor2_2 _10423_ (.A(_04538_),
    .B(_04541_),
    .Y(_04590_));
 sky130_fd_sc_hd__xnor2_1 _10424_ (.A(_04533_),
    .B(_04536_),
    .Y(_04591_));
 sky130_fd_sc_hd__xor2_2 _10425_ (.A(_04375_),
    .B(_04531_),
    .X(_04592_));
 sky130_fd_sc_hd__inv_2 _10426_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__xnor2_2 _10427_ (.A(_04525_),
    .B(_04528_),
    .Y(_04594_));
 sky130_fd_sc_hd__inv_2 _10428_ (.A(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__xnor2_2 _10429_ (.A(_04520_),
    .B(_04524_),
    .Y(_04596_));
 sky130_fd_sc_hd__inv_2 _10430_ (.A(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__xnor2_1 _10431_ (.A(_04515_),
    .B(_04518_),
    .Y(_04599_));
 sky130_fd_sc_hd__inv_2 _10432_ (.A(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__xor2_1 _10433_ (.A(_04395_),
    .B(_04514_),
    .X(_04601_));
 sky130_fd_sc_hd__xnor2_1 _10434_ (.A(_04395_),
    .B(_04514_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _10435_ (.A(_04398_),
    .B(_04399_),
    .Y(_04603_));
 sky130_fd_sc_hd__xnor2_2 _10436_ (.A(_04512_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__xnor2_2 _10437_ (.A(_04403_),
    .B(_04509_),
    .Y(_04605_));
 sky130_fd_sc_hd__inv_2 _10438_ (.A(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_1 _10439_ (.A(_04407_),
    .B(_04408_),
    .Y(_04607_));
 sky130_fd_sc_hd__xor2_2 _10440_ (.A(_04507_),
    .B(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__nor2_1 _10441_ (.A(_04415_),
    .B(_04417_),
    .Y(_04610_));
 sky130_fd_sc_hd__xnor2_2 _10442_ (.A(_04505_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _10443_ (.A(_04425_),
    .B(_04426_),
    .Y(_04612_));
 sky130_fd_sc_hd__xor2_2 _10444_ (.A(_04503_),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__xnor2_2 _10445_ (.A(_04497_),
    .B(_04500_),
    .Y(_04614_));
 sky130_fd_sc_hd__and3_1 _10446_ (.A(_04494_),
    .B(_04457_),
    .C(_04456_),
    .X(_04615_));
 sky130_fd_sc_hd__a21oi_2 _10447_ (.A1(_04456_),
    .A2(_04457_),
    .B1(_04494_),
    .Y(_04616_));
 sky130_fd_sc_hd__nor2_1 _10448_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__a22o_1 _10449_ (.A1(_04464_),
    .A2(_04465_),
    .B1(_04474_),
    .B2(_04492_),
    .X(_04618_));
 sky130_fd_sc_hd__and2_1 _10450_ (.A(_04493_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_04474_),
    .B(_04475_),
    .Y(_04621_));
 sky130_fd_sc_hd__xnor2_2 _10452_ (.A(_04491_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__or4b_1 _10453_ (.A(_04575_),
    .B(_04580_),
    .C(_04619_),
    .D_N(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__a21oi_1 _10454_ (.A1(_04456_),
    .A2(_04495_),
    .B1(_04450_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor2_1 _10455_ (.A(_04496_),
    .B(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_04430_),
    .B(_04431_),
    .Y(_04626_));
 sky130_fd_sc_hd__xnor2_2 _10457_ (.A(_04501_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__nor4b_1 _10458_ (.A(_04611_),
    .B(_04613_),
    .C(_04625_),
    .D_N(_04617_),
    .Y(_04628_));
 sky130_fd_sc_hd__and4bb_1 _10459_ (.A_N(_04623_),
    .B_N(_04627_),
    .C(_04614_),
    .D(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__or4bb_1 _10460_ (.A(_04604_),
    .B(_04605_),
    .C_N(_04608_),
    .D_N(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__or4_1 _10461_ (.A(_04600_),
    .B(_04630_),
    .C(_04601_),
    .D(_04597_),
    .X(_04632_));
 sky130_fd_sc_hd__and4b_1 _10462_ (.A_N(_04632_),
    .B(_04594_),
    .C(_04592_),
    .D(_04591_),
    .X(_04633_));
 sky130_fd_sc_hd__nand3_1 _10463_ (.A(_04585_),
    .B(_04590_),
    .C(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__a211oi_4 _10464_ (.A1(_04561_),
    .A2(_04586_),
    .B1(_04589_),
    .C1(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand3_4 _10465_ (.A(net100),
    .B(_04583_),
    .C(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o31ai_1 _10466_ (.A1(_00803_),
    .A2(_00891_),
    .A3(_03618_),
    .B1(_00748_),
    .Y(_04637_));
 sky130_fd_sc_hd__a31oi_1 _10467_ (.A1(_04584_),
    .A2(_04636_),
    .A3(_03601_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__o32ai_2 _10468_ (.A1(_03606_),
    .A2(_03614_),
    .A3(_03611_),
    .B1(net65),
    .B2(_04638_),
    .Y(net67));
 sky130_fd_sc_hd__and4_1 _10469_ (.A(_03552_),
    .B(_01694_),
    .C(_01958_),
    .D(_03613_),
    .X(_04639_));
 sky130_fd_sc_hd__xnor2_4 _10470_ (.A(_03512_),
    .B(_03514_),
    .Y(_04640_));
 sky130_fd_sc_hd__a211o_1 _10471_ (.A1(_03554_),
    .A2(_04640_),
    .B1(_04639_),
    .C1(net103),
    .X(_04642_));
 sky130_fd_sc_hd__and3_4 _10472_ (.A(_03601_),
    .B(_05339_),
    .C(_00748_),
    .X(_04643_));
 sky130_fd_sc_hd__or3_2 _10473_ (.A(net65),
    .B(_00517_),
    .C(_00638_),
    .X(_04644_));
 sky130_fd_sc_hd__a31o_4 _10474_ (.A1(net100),
    .A2(_04583_),
    .A3(_04635_),
    .B1(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__a21oi_1 _10475_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04581_),
    .Y(_04646_));
 sky130_fd_sc_hd__a311o_1 _10476_ (.A1(_04568_),
    .A2(_04575_),
    .A3(_04582_),
    .B1(_04646_),
    .C1(_04572_),
    .X(_04647_));
 sky130_fd_sc_hd__a21oi_1 _10477_ (.A1(_04572_),
    .A2(_04622_),
    .B1(_04645_),
    .Y(_04648_));
 sky130_fd_sc_hd__a2bb2o_1 _10478_ (.A1_N(net99),
    .A2_N(_04642_),
    .B1(_04647_),
    .B2(_04648_),
    .X(net78));
 sky130_fd_sc_hd__and4_1 _10479_ (.A(_03552_),
    .B(_01694_),
    .C(_01958_),
    .D(_04640_),
    .X(_04649_));
 sky130_fd_sc_hd__xnor2_4 _10480_ (.A(_01493_),
    .B(_03515_),
    .Y(_04650_));
 sky130_fd_sc_hd__a211o_1 _10481_ (.A1(_03554_),
    .A2(_04650_),
    .B1(_04649_),
    .C1(net103),
    .X(_04652_));
 sky130_fd_sc_hd__a21o_1 _10482_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04577_),
    .X(_04653_));
 sky130_fd_sc_hd__o211a_1 _10483_ (.A1(_04622_),
    .A2(_04583_),
    .B1(_04573_),
    .C1(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__a21oi_2 _10484_ (.A1(_04493_),
    .A2(_04618_),
    .B1(_04573_),
    .Y(_04655_));
 sky130_fd_sc_hd__o32ai_4 _10485_ (.A1(_04655_),
    .A2(_04645_),
    .A3(_04654_),
    .B1(_04652_),
    .B2(net99),
    .Y(net89));
 sky130_fd_sc_hd__nand2_2 _10486_ (.A(_01308_),
    .B(_01310_),
    .Y(_04656_));
 sky130_fd_sc_hd__xnor2_4 _10487_ (.A(_03517_),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _10488_ (.A(_03554_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__o211a_1 _10489_ (.A1(_03554_),
    .A2(_04650_),
    .B1(_04658_),
    .C1(_03612_),
    .X(_04659_));
 sky130_fd_sc_hd__nand2_1 _10490_ (.A(_04583_),
    .B(_04622_),
    .Y(_04660_));
 sky130_fd_sc_hd__o21ai_1 _10491_ (.A1(_04583_),
    .A2(_04619_),
    .B1(_04660_),
    .Y(_04662_));
 sky130_fd_sc_hd__o211a_1 _10492_ (.A1(_03618_),
    .A2(_04570_),
    .B1(_04617_),
    .C1(_04569_),
    .X(_04663_));
 sky130_fd_sc_hd__a211o_1 _10493_ (.A1(_04662_),
    .A2(_04573_),
    .B1(_04663_),
    .C1(_04645_),
    .X(_04664_));
 sky130_fd_sc_hd__o31ai_2 _10494_ (.A1(net103),
    .A2(_04659_),
    .A3(net99),
    .B1(_04664_),
    .Y(net92));
 sky130_fd_sc_hd__o211a_1 _10495_ (.A1(_04615_),
    .A2(_04616_),
    .B1(_04568_),
    .C1(_04582_),
    .X(_04665_));
 sky130_fd_sc_hd__a211o_1 _10496_ (.A1(_04619_),
    .A2(_04583_),
    .B1(_04572_),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__o2111ai_2 _10497_ (.A1(_04573_),
    .A2(_04625_),
    .B1(_04636_),
    .C1(_04643_),
    .D1(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__a21o_1 _10498_ (.A1(_01308_),
    .A2(_03518_),
    .B1(_01124_),
    .X(_04668_));
 sky130_fd_sc_hd__nand2_4 _10499_ (.A(_03519_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _10500_ (.A(_03555_),
    .B(_04657_),
    .Y(_04670_));
 sky130_fd_sc_hd__o211a_1 _10501_ (.A1(_04669_),
    .A2(_03555_),
    .B1(_03612_),
    .C1(_04670_),
    .X(_04672_));
 sky130_fd_sc_hd__o31ai_2 _10502_ (.A1(net103),
    .A2(_04672_),
    .A3(net99),
    .B1(_04667_),
    .Y(net93));
 sky130_fd_sc_hd__nor2_1 _10503_ (.A(_04573_),
    .B(_04614_),
    .Y(_04673_));
 sky130_fd_sc_hd__a211o_1 _10504_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04615_),
    .C1(_04616_),
    .X(_04674_));
 sky130_fd_sc_hd__o211a_1 _10505_ (.A1(_04625_),
    .A2(_04583_),
    .B1(_04573_),
    .C1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__o21bai_1 _10506_ (.A1(_04673_),
    .A2(_04675_),
    .B1_N(_04645_),
    .Y(_04676_));
 sky130_fd_sc_hd__xor2_4 _10507_ (.A(_03521_),
    .B(_03523_),
    .X(_04677_));
 sky130_fd_sc_hd__a31o_1 _10508_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__o211a_1 _10509_ (.A1(_03554_),
    .A2(_04669_),
    .B1(_04678_),
    .C1(_03612_),
    .X(_04679_));
 sky130_fd_sc_hd__o31ai_2 _10510_ (.A1(net103),
    .A2(_04679_),
    .A3(net99),
    .B1(_04676_),
    .Y(net94));
 sky130_fd_sc_hd__a211o_1 _10511_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04624_),
    .C1(_04496_),
    .X(_04681_));
 sky130_fd_sc_hd__nor2_1 _10512_ (.A(_04573_),
    .B(_04627_),
    .Y(_04682_));
 sky130_fd_sc_hd__o211a_1 _10513_ (.A1(_04583_),
    .A2(_04614_),
    .B1(_04681_),
    .C1(_04573_),
    .X(_04683_));
 sky130_fd_sc_hd__xnor2_4 _10514_ (.A(_00740_),
    .B(_03524_),
    .Y(_04684_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(_04677_),
    .A1(_04684_),
    .S(_03554_),
    .X(_04685_));
 sky130_fd_sc_hd__or2_1 _10516_ (.A(net103),
    .B(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__o32ai_4 _10517_ (.A1(_04645_),
    .A2(_04682_),
    .A3(_04683_),
    .B1(_04686_),
    .B2(net99),
    .Y(net95));
 sky130_fd_sc_hd__xor2_4 _10518_ (.A(_03525_),
    .B(_03527_),
    .X(_04687_));
 sky130_fd_sc_hd__a31o_1 _10519_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__o211a_1 _10520_ (.A1(_03554_),
    .A2(_04684_),
    .B1(_04688_),
    .C1(_03612_),
    .X(_04689_));
 sky130_fd_sc_hd__nand2_1 _10521_ (.A(_04583_),
    .B(_04614_),
    .Y(_04691_));
 sky130_fd_sc_hd__o211a_1 _10522_ (.A1(_04583_),
    .A2(_04627_),
    .B1(_04691_),
    .C1(_04573_),
    .X(_04692_));
 sky130_fd_sc_hd__a21oi_1 _10523_ (.A1(_04572_),
    .A2(_04613_),
    .B1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__o32ai_4 _10524_ (.A1(net103),
    .A2(_04689_),
    .A3(net99),
    .B1(_04693_),
    .B2(_04645_),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_2 _10525_ (.A(_00411_),
    .B(_03528_),
    .Y(_04694_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(_04687_),
    .A1(_04694_),
    .S(_03554_),
    .X(_04695_));
 sky130_fd_sc_hd__a21o_1 _10527_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04627_),
    .X(_04696_));
 sky130_fd_sc_hd__nand2_1 _10528_ (.A(_04572_),
    .B(_04611_),
    .Y(_04697_));
 sky130_fd_sc_hd__o211ai_1 _10529_ (.A1(_04583_),
    .A2(_04613_),
    .B1(_04696_),
    .C1(_04573_),
    .Y(_04698_));
 sky130_fd_sc_hd__a21o_1 _10530_ (.A1(_04697_),
    .A2(_04698_),
    .B1(_04645_),
    .X(_04699_));
 sky130_fd_sc_hd__o31ai_2 _10531_ (.A1(net103),
    .A2(_04695_),
    .A3(net99),
    .B1(_04699_),
    .Y(net97));
 sky130_fd_sc_hd__xnor2_2 _10532_ (.A(_03529_),
    .B(_03530_),
    .Y(_04701_));
 sky130_fd_sc_hd__a31o_1 _10533_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__o211a_1 _10534_ (.A1(_03554_),
    .A2(_04694_),
    .B1(_04702_),
    .C1(_03612_),
    .X(_04703_));
 sky130_fd_sc_hd__nand3_1 _10535_ (.A(_04568_),
    .B(_04582_),
    .C(_04611_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21boi_1 _10536_ (.A1(_04583_),
    .A2(_04613_),
    .B1_N(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__o211a_1 _10537_ (.A1(_03618_),
    .A2(_04570_),
    .B1(_04608_),
    .C1(_04569_),
    .X(_04706_));
 sky130_fd_sc_hd__a211o_1 _10538_ (.A1(_04573_),
    .A2(_04705_),
    .B1(_04706_),
    .C1(_04645_),
    .X(_04707_));
 sky130_fd_sc_hd__o31ai_2 _10539_ (.A1(net104),
    .A2(_04703_),
    .A3(net99),
    .B1(_04707_),
    .Y(net98));
 sky130_fd_sc_hd__a221o_1 _10540_ (.A1(_03617_),
    .A2(_04571_),
    .B1(_04568_),
    .B2(_04347_),
    .C1(_04606_),
    .X(_04708_));
 sky130_fd_sc_hd__nand2_1 _10541_ (.A(_04583_),
    .B(_04611_),
    .Y(_04710_));
 sky130_fd_sc_hd__o21a_1 _10542_ (.A1(_04583_),
    .A2(_04608_),
    .B1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__o21a_1 _10543_ (.A1(_04572_),
    .A2(_04711_),
    .B1(_04708_),
    .X(_04712_));
 sky130_fd_sc_hd__xnor2_2 _10544_ (.A(_00141_),
    .B(_03532_),
    .Y(_04713_));
 sky130_fd_sc_hd__a31o_1 _10545_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__o211a_1 _10546_ (.A1(_03554_),
    .A2(_04701_),
    .B1(_04714_),
    .C1(_03612_),
    .X(_04715_));
 sky130_fd_sc_hd__o32ai_4 _10547_ (.A1(net104),
    .A2(_04715_),
    .A3(net99),
    .B1(_04645_),
    .B2(_04712_),
    .Y(net68));
 sky130_fd_sc_hd__o211a_1 _10548_ (.A1(_03618_),
    .A2(_04570_),
    .B1(_04604_),
    .C1(_04569_),
    .X(_04716_));
 sky130_fd_sc_hd__a21oi_1 _10549_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04608_),
    .Y(_04717_));
 sky130_fd_sc_hd__a31o_1 _10550_ (.A1(_04568_),
    .A2(_04582_),
    .A3(_04605_),
    .B1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a21oi_2 _10551_ (.A1(_04573_),
    .A2(_04718_),
    .B1(_04716_),
    .Y(_04720_));
 sky130_fd_sc_hd__a21oi_1 _10552_ (.A1(_00031_),
    .A2(_00032_),
    .B1(_03533_),
    .Y(_04721_));
 sky130_fd_sc_hd__and3_1 _10553_ (.A(_03533_),
    .B(_00032_),
    .C(_00031_),
    .X(_04722_));
 sky130_fd_sc_hd__nor2_1 _10554_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__a31o_1 _10555_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__o211a_1 _10556_ (.A1(_03554_),
    .A2(_04713_),
    .B1(_04724_),
    .C1(_03612_),
    .X(_04725_));
 sky130_fd_sc_hd__o32ai_4 _10557_ (.A1(net104),
    .A2(_04725_),
    .A3(net99),
    .B1(_04645_),
    .B2(_04720_),
    .Y(net69));
 sky130_fd_sc_hd__nand3_1 _10558_ (.A(_04568_),
    .B(_04582_),
    .C(_04604_),
    .Y(_04726_));
 sky130_fd_sc_hd__a21boi_1 _10559_ (.A1(_04583_),
    .A2(_04605_),
    .B1_N(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(_04727_),
    .A1(_04602_),
    .S(_04572_),
    .X(_04728_));
 sky130_fd_sc_hd__xor2_2 _10561_ (.A(_05274_),
    .B(_03535_),
    .X(_04730_));
 sky130_fd_sc_hd__a31o_1 _10562_ (.A1(_03552_),
    .A2(_01694_),
    .A3(_01958_),
    .B1(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__o211a_1 _10563_ (.A1(_04723_),
    .A2(_03554_),
    .B1(_03612_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__o32ai_4 _10564_ (.A1(net104),
    .A2(_04732_),
    .A3(net99),
    .B1(_04645_),
    .B2(_04728_),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_2 _10565_ (.A(_03536_),
    .B(_03538_),
    .Y(_04733_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(_04730_),
    .A1(_04733_),
    .S(_03554_),
    .X(_04734_));
 sky130_fd_sc_hd__a21o_1 _10567_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04604_),
    .X(_04735_));
 sky130_fd_sc_hd__o211a_1 _10568_ (.A1(_04601_),
    .A2(_04583_),
    .B1(net100),
    .C1(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__a21oi_1 _10569_ (.A1(_04572_),
    .A2(_04600_),
    .B1(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__o32ai_4 _10570_ (.A1(net105),
    .A2(_04734_),
    .A3(net99),
    .B1(_04737_),
    .B2(_04645_),
    .Y(net71));
 sky130_fd_sc_hd__nand3_1 _10571_ (.A(_04568_),
    .B(_04582_),
    .C(_04600_),
    .Y(_04739_));
 sky130_fd_sc_hd__a21boi_1 _10572_ (.A1(_04583_),
    .A2(_04601_),
    .B1_N(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(_04740_),
    .A1(_04596_),
    .S(_04572_),
    .X(_04741_));
 sky130_fd_sc_hd__xnor2_1 _10574_ (.A(_05096_),
    .B(_03539_),
    .Y(_04742_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(_04733_),
    .A1(_04742_),
    .S(_03554_),
    .X(_04743_));
 sky130_fd_sc_hd__or2_1 _10576_ (.A(net104),
    .B(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__o22ai_2 _10577_ (.A1(net99),
    .A2(_04744_),
    .B1(_04645_),
    .B2(_04741_),
    .Y(net72));
 sky130_fd_sc_hd__a21boi_1 _10578_ (.A1(_03539_),
    .A2(_05096_),
    .B1_N(_05095_),
    .Y(_04745_));
 sky130_fd_sc_hd__xnor2_2 _10579_ (.A(_05013_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__nor2_1 _10580_ (.A(_04746_),
    .B(_03555_),
    .Y(_04747_));
 sky130_fd_sc_hd__and4_1 _10581_ (.A(_03552_),
    .B(_01694_),
    .C(_01958_),
    .D(_04742_),
    .X(_04749_));
 sky130_fd_sc_hd__a21o_1 _10582_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04599_),
    .X(_04750_));
 sky130_fd_sc_hd__o211a_1 _10583_ (.A1(_04583_),
    .A2(_04596_),
    .B1(_04750_),
    .C1(net100),
    .X(_04751_));
 sky130_fd_sc_hd__a211o_1 _10584_ (.A1(_04572_),
    .A2(_04594_),
    .B1(_04645_),
    .C1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__o41ai_2 _10585_ (.A1(net105),
    .A2(_04747_),
    .A3(_04749_),
    .A4(net99),
    .B1(_04752_),
    .Y(net73));
 sky130_fd_sc_hd__xnor2_1 _10586_ (.A(_03541_),
    .B(_03543_),
    .Y(_04753_));
 sky130_fd_sc_hd__nor2_1 _10587_ (.A(_03554_),
    .B(_04746_),
    .Y(_04754_));
 sky130_fd_sc_hd__a211o_1 _10588_ (.A1(_03554_),
    .A2(_04753_),
    .B1(_04754_),
    .C1(net105),
    .X(_04755_));
 sky130_fd_sc_hd__a21o_1 _10589_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04597_),
    .X(_04756_));
 sky130_fd_sc_hd__o211a_1 _10590_ (.A1(_04595_),
    .A2(_04583_),
    .B1(net100),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a21oi_1 _10591_ (.A1(_04572_),
    .A2(_04593_),
    .B1(_04757_),
    .Y(_04759_));
 sky130_fd_sc_hd__o22ai_2 _10592_ (.A1(net99),
    .A2(_04755_),
    .B1(_04759_),
    .B2(_04645_),
    .Y(net74));
 sky130_fd_sc_hd__xor2_1 _10593_ (.A(_04777_),
    .B(_03544_),
    .X(_04760_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(_04753_),
    .A1(_04760_),
    .S(_03554_),
    .X(_04761_));
 sky130_fd_sc_hd__a21o_1 _10595_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04595_),
    .X(_04762_));
 sky130_fd_sc_hd__o211ai_1 _10596_ (.A1(_04593_),
    .A2(_04583_),
    .B1(net100),
    .C1(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__o21a_1 _10597_ (.A1(net100),
    .A2(_04591_),
    .B1(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__o32ai_4 _10598_ (.A1(net105),
    .A2(_04761_),
    .A3(_03606_),
    .B1(_04764_),
    .B2(_04645_),
    .Y(net75));
 sky130_fd_sc_hd__xnor2_1 _10599_ (.A(_04180_),
    .B(_03545_),
    .Y(_04765_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(_04760_),
    .A1(_04765_),
    .S(_03554_),
    .X(_04766_));
 sky130_fd_sc_hd__and3_1 _10601_ (.A(_04568_),
    .B(_04582_),
    .C(_04591_),
    .X(_04768_));
 sky130_fd_sc_hd__a21oi_1 _10602_ (.A1(_04583_),
    .A2(_04592_),
    .B1(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _10603_ (.A(_04572_),
    .B(_04590_),
    .Y(_04770_));
 sky130_fd_sc_hd__o21ai_1 _10604_ (.A1(_04572_),
    .A2(_04769_),
    .B1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__o32ai_4 _10605_ (.A1(net105),
    .A2(_04766_),
    .A3(_03606_),
    .B1(_04771_),
    .B2(_04645_),
    .Y(net76));
 sky130_fd_sc_hd__xor2_1 _10606_ (.A(_03586_),
    .B(_03546_),
    .X(_04772_));
 sky130_fd_sc_hd__inv_2 _10607_ (.A(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(_04765_),
    .A1(_04773_),
    .S(_03554_),
    .X(_04774_));
 sky130_fd_sc_hd__a21o_1 _10609_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04591_),
    .X(_04775_));
 sky130_fd_sc_hd__o21ai_1 _10610_ (.A1(_04583_),
    .A2(_04590_),
    .B1(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(_04572_),
    .B(_04585_),
    .Y(_04778_));
 sky130_fd_sc_hd__o21ai_1 _10612_ (.A1(_04572_),
    .A2(_04776_),
    .B1(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__o32ai_2 _10613_ (.A1(_03606_),
    .A2(_04774_),
    .A3(_03611_),
    .B1(_04645_),
    .B2(_04779_),
    .Y(net77));
 sky130_fd_sc_hd__xor2_1 _10614_ (.A(_03047_),
    .B(_03547_),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(_04773_),
    .A1(_04780_),
    .S(_03554_),
    .X(_04781_));
 sky130_fd_sc_hd__a21o_1 _10616_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04590_),
    .X(_04782_));
 sky130_fd_sc_hd__o211ai_1 _10617_ (.A1(_04583_),
    .A2(_04585_),
    .B1(_04782_),
    .C1(net100),
    .Y(_04783_));
 sky130_fd_sc_hd__o21ai_1 _10618_ (.A1(net100),
    .A2(_04589_),
    .B1(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__o32ai_2 _10619_ (.A1(_03611_),
    .A2(_04781_),
    .A3(_03606_),
    .B1(_04784_),
    .B2(_04645_),
    .Y(net79));
 sky130_fd_sc_hd__xnor2_1 _10620_ (.A(_02552_),
    .B(_03548_),
    .Y(_04785_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(_04780_),
    .A1(_04785_),
    .S(_03554_),
    .X(_04787_));
 sky130_fd_sc_hd__a21o_1 _10622_ (.A1(_04561_),
    .A2(_04586_),
    .B1(net100),
    .X(_04788_));
 sky130_fd_sc_hd__nand3_1 _10623_ (.A(net100),
    .B(_04583_),
    .C(_04585_),
    .Y(_04789_));
 sky130_fd_sc_hd__o311ai_2 _10624_ (.A1(_04572_),
    .A2(_04589_),
    .A3(_04583_),
    .B1(_04789_),
    .C1(_04788_),
    .Y(_04790_));
 sky130_fd_sc_hd__o32ai_2 _10625_ (.A1(_03611_),
    .A2(_04787_),
    .A3(_03606_),
    .B1(_04790_),
    .B2(_04645_),
    .Y(net80));
 sky130_fd_sc_hd__a2111o_1 _10626_ (.A1(_03548_),
    .A2(_02552_),
    .B1(_02530_),
    .C1(_03551_),
    .D1(_03550_),
    .X(_04791_));
 sky130_fd_sc_hd__a21boi_1 _10627_ (.A1(_03552_),
    .A2(_04791_),
    .B1_N(_03554_),
    .Y(_04792_));
 sky130_fd_sc_hd__a211oi_1 _10628_ (.A1(_04785_),
    .A2(_03555_),
    .B1(_03611_),
    .C1(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__a41oi_2 _10629_ (.A1(_03598_),
    .A2(_03600_),
    .A3(_03601_),
    .A4(_04793_),
    .B1(_00924_),
    .Y(_04794_));
 sky130_fd_sc_hd__a211oi_1 _10630_ (.A1(_04561_),
    .A2(_04586_),
    .B1(_04583_),
    .C1(_04572_),
    .Y(_04795_));
 sky130_fd_sc_hd__o31a_1 _10631_ (.A1(_04555_),
    .A2(_04572_),
    .A3(_04588_),
    .B1(_04583_),
    .X(_04797_));
 sky130_fd_sc_hd__o32ai_2 _10632_ (.A1(_04644_),
    .A2(_04795_),
    .A3(_04797_),
    .B1(_05339_),
    .B2(_04794_),
    .Y(net81));
 sky130_fd_sc_hd__nand3_1 _10633_ (.A(_03557_),
    .B(_03577_),
    .C(_03612_),
    .Y(_04798_));
 sky130_fd_sc_hd__a21oi_1 _10634_ (.A1(_03598_),
    .A2(_04798_),
    .B1(_03599_),
    .Y(_04799_));
 sky130_fd_sc_hd__mux2_4 _10635_ (.A0(net16),
    .A1(net48),
    .S(_03651_),
    .X(_04800_));
 sky130_fd_sc_hd__nand4_1 _10636_ (.A(net100),
    .B(_04800_),
    .C(_04582_),
    .D(_04568_),
    .Y(_04801_));
 sky130_fd_sc_hd__o21bai_1 _10637_ (.A1(_04583_),
    .A2(_04572_),
    .B1_N(_04800_),
    .Y(_04802_));
 sky130_fd_sc_hd__a32o_1 _10638_ (.A1(net100),
    .A2(_04635_),
    .A3(_04583_),
    .B1(_04802_),
    .B2(_04801_),
    .X(_04803_));
 sky130_fd_sc_hd__a2bb2oi_1 _10639_ (.A1_N(_03604_),
    .A2_N(_04799_),
    .B1(_04803_),
    .B2(_04643_),
    .Y(net82));
 sky130_fd_sc_hd__a21oi_1 _10640_ (.A1(_03557_),
    .A2(_03558_),
    .B1(_03611_),
    .Y(_04804_));
 sky130_fd_sc_hd__o21ai_1 _10641_ (.A1(_03557_),
    .A2(_03558_),
    .B1(_04804_),
    .Y(_04806_));
 sky130_fd_sc_hd__a21o_1 _10642_ (.A1(_03598_),
    .A2(_04806_),
    .B1(_03599_),
    .X(_04807_));
 sky130_fd_sc_hd__mux2_2 _10643_ (.A0(net17),
    .A1(net49),
    .S(_03651_),
    .X(_04808_));
 sky130_fd_sc_hd__nand3_1 _10644_ (.A(_04568_),
    .B(_04582_),
    .C(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_1 _10645_ (.A(_04800_),
    .B(_04808_),
    .Y(_04810_));
 sky130_fd_sc_hd__and2_1 _10646_ (.A(_04800_),
    .B(_04808_),
    .X(_04811_));
 sky130_fd_sc_hd__nor2_1 _10647_ (.A(_04810_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _10648_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__a21oi_1 _10649_ (.A1(_04635_),
    .A2(_04583_),
    .B1(_04572_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand3_1 _10650_ (.A(net100),
    .B(_04809_),
    .C(_04813_),
    .Y(_04815_));
 sky130_fd_sc_hd__o211ai_1 _10651_ (.A1(_04812_),
    .A2(net100),
    .B1(_04636_),
    .C1(_04815_),
    .Y(_04817_));
 sky130_fd_sc_hd__a22oi_1 _10652_ (.A1(_04817_),
    .A2(_04643_),
    .B1(_04807_),
    .B2(_03603_),
    .Y(net83));
 sky130_fd_sc_hd__a221o_1 _10653_ (.A1(_03556_),
    .A2(_03559_),
    .B1(_03561_),
    .B2(_03590_),
    .C1(_03611_),
    .X(_04818_));
 sky130_fd_sc_hd__a21o_1 _10654_ (.A1(_03598_),
    .A2(_04818_),
    .B1(_03599_),
    .X(_04819_));
 sky130_fd_sc_hd__mux2_4 _10655_ (.A0(net18),
    .A1(net50),
    .S(_03651_),
    .X(_04820_));
 sky130_fd_sc_hd__nor3_1 _10656_ (.A(_04800_),
    .B(_04808_),
    .C(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21boi_1 _10657_ (.A1(_04583_),
    .A2(_04810_),
    .B1_N(_04820_),
    .Y(_04822_));
 sky130_fd_sc_hd__xor2_1 _10658_ (.A(_04811_),
    .B(_04820_),
    .X(_04823_));
 sky130_fd_sc_hd__a21o_1 _10659_ (.A1(_04583_),
    .A2(_04821_),
    .B1(_04572_),
    .X(_04824_));
 sky130_fd_sc_hd__o221ai_1 _10660_ (.A1(net100),
    .A2(_04823_),
    .B1(_04822_),
    .B2(_04824_),
    .C1(_04636_),
    .Y(_04825_));
 sky130_fd_sc_hd__a22oi_1 _10661_ (.A1(_04825_),
    .A2(_04643_),
    .B1(_04819_),
    .B2(_03603_),
    .Y(net84));
 sky130_fd_sc_hd__nand3_1 _10662_ (.A(_03566_),
    .B(_03591_),
    .C(_03612_),
    .Y(_04827_));
 sky130_fd_sc_hd__a21o_1 _10663_ (.A1(_03598_),
    .A2(_04827_),
    .B1(_03599_),
    .X(_04828_));
 sky130_fd_sc_hd__mux2_2 _10664_ (.A0(net19),
    .A1(net51),
    .S(_03651_),
    .X(_04829_));
 sky130_fd_sc_hd__nor4_4 _10665_ (.A(_04800_),
    .B(_04808_),
    .C(_04820_),
    .D(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__inv_2 _10666_ (.A(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__a21oi_1 _10667_ (.A1(_04568_),
    .A2(_04582_),
    .B1(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21o_1 _10668_ (.A1(_04583_),
    .A2(_04830_),
    .B1(_04572_),
    .X(_04833_));
 sky130_fd_sc_hd__a21boi_1 _10669_ (.A1(_04583_),
    .A2(_04821_),
    .B1_N(_04829_),
    .Y(_04834_));
 sky130_fd_sc_hd__a21oi_1 _10670_ (.A1(_04811_),
    .A2(_04820_),
    .B1(_04829_),
    .Y(_04835_));
 sky130_fd_sc_hd__and3_1 _10671_ (.A(_04811_),
    .B(_04820_),
    .C(_04829_),
    .X(_04837_));
 sky130_fd_sc_hd__o21ai_1 _10672_ (.A1(_04835_),
    .A2(_04837_),
    .B1(_04572_),
    .Y(_04838_));
 sky130_fd_sc_hd__o211ai_1 _10673_ (.A1(_04834_),
    .A2(_04833_),
    .B1(_04636_),
    .C1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__a22oi_1 _10674_ (.A1(_04839_),
    .A2(_04643_),
    .B1(_04828_),
    .B2(_03603_),
    .Y(net85));
 sky130_fd_sc_hd__nand3_1 _10675_ (.A(_03568_),
    .B(_03576_),
    .C(_03612_),
    .Y(_04840_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(_03598_),
    .A2(_04840_),
    .B1(_03599_),
    .X(_04841_));
 sky130_fd_sc_hd__a311o_1 _10677_ (.A1(_03633_),
    .A2(_03635_),
    .A3(_03637_),
    .B1(net115),
    .C1(net52),
    .X(_04842_));
 sky130_fd_sc_hd__o21a_1 _10678_ (.A1(net20),
    .A2(_03651_),
    .B1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__o21ai_2 _10679_ (.A1(net20),
    .A2(_03651_),
    .B1(_04842_),
    .Y(_04844_));
 sky130_fd_sc_hd__a31o_1 _10680_ (.A1(_04811_),
    .A2(_04820_),
    .A3(_04829_),
    .B1(_04843_),
    .X(_04845_));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_04837_),
    .B(_04843_),
    .Y(_04847_));
 sky130_fd_sc_hd__a21o_1 _10682_ (.A1(_04845_),
    .A2(_04847_),
    .B1(net100),
    .X(_04848_));
 sky130_fd_sc_hd__a21oi_1 _10683_ (.A1(_04583_),
    .A2(_04830_),
    .B1(_04844_),
    .Y(_04849_));
 sky130_fd_sc_hd__a31o_1 _10684_ (.A1(_04583_),
    .A2(_04830_),
    .A3(_04844_),
    .B1(_04572_),
    .X(_04850_));
 sky130_fd_sc_hd__o211ai_1 _10685_ (.A1(_04849_),
    .A2(_04850_),
    .B1(_04636_),
    .C1(_04848_),
    .Y(_04851_));
 sky130_fd_sc_hd__a22oi_1 _10686_ (.A1(_04851_),
    .A2(_04643_),
    .B1(_03603_),
    .B2(_04841_),
    .Y(net86));
 sky130_fd_sc_hd__o211ai_1 _10687_ (.A1(_01364_),
    .A2(_03566_),
    .B1(_03594_),
    .C1(_03612_),
    .Y(_04852_));
 sky130_fd_sc_hd__a21o_1 _10688_ (.A1(_03598_),
    .A2(_04852_),
    .B1(_03599_),
    .X(_04853_));
 sky130_fd_sc_hd__a21oi_1 _10689_ (.A1(_03643_),
    .A2(_03649_),
    .B1(net21),
    .Y(_04854_));
 sky130_fd_sc_hd__o311a_1 _10690_ (.A1(_03636_),
    .A2(_03638_),
    .A3(_03632_),
    .B1(_03649_),
    .C1(_00286_),
    .X(_04855_));
 sky130_fd_sc_hd__a21oi_1 _10691_ (.A1(_00286_),
    .A2(_03651_),
    .B1(_04854_),
    .Y(_04857_));
 sky130_fd_sc_hd__o21a_1 _10692_ (.A1(_04854_),
    .A2(_04855_),
    .B1(_04844_),
    .X(_04858_));
 sky130_fd_sc_hd__and3_1 _10693_ (.A(_04583_),
    .B(_04830_),
    .C(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__a21boi_1 _10694_ (.A1(_04832_),
    .A2(_04844_),
    .B1_N(_04857_),
    .Y(_04860_));
 sky130_fd_sc_hd__o21ai_1 _10695_ (.A1(_04859_),
    .A2(_04860_),
    .B1(_04814_),
    .Y(_04861_));
 sky130_fd_sc_hd__and3_1 _10696_ (.A(_04837_),
    .B(_04843_),
    .C(_04857_),
    .X(_04862_));
 sky130_fd_sc_hd__o2bb2a_1 _10697_ (.A1_N(_04837_),
    .A2_N(_04843_),
    .B1(_04854_),
    .B2(_04855_),
    .X(_04863_));
 sky130_fd_sc_hd__o31a_1 _10698_ (.A1(_04862_),
    .A2(_04863_),
    .A3(net100),
    .B1(_04643_),
    .X(_04864_));
 sky130_fd_sc_hd__a22oi_1 _10699_ (.A1(_04861_),
    .A2(_04864_),
    .B1(_04853_),
    .B2(_03603_),
    .Y(net87));
 sky130_fd_sc_hd__and3_1 _10700_ (.A(_03573_),
    .B(_03574_),
    .C(_03600_),
    .X(_04865_));
 sky130_fd_sc_hd__o21ai_1 _10701_ (.A1(_03612_),
    .A2(_03595_),
    .B1(_04865_),
    .Y(_04867_));
 sky130_fd_sc_hd__a311o_1 _10702_ (.A1(_03633_),
    .A2(_03635_),
    .A3(_03637_),
    .B1(net115),
    .C1(net54),
    .X(_04868_));
 sky130_fd_sc_hd__o21a_1 _10703_ (.A1(net22),
    .A2(_03651_),
    .B1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__o21ai_2 _10704_ (.A1(net22),
    .A2(_03651_),
    .B1(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__and4_1 _10705_ (.A(_04583_),
    .B(_04830_),
    .C(_04858_),
    .D(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a21oi_1 _10706_ (.A1(_04832_),
    .A2(_04858_),
    .B1(_04870_),
    .Y(_04872_));
 sky130_fd_sc_hd__o21ai_1 _10707_ (.A1(_04871_),
    .A2(_04872_),
    .B1(_04814_),
    .Y(_04873_));
 sky130_fd_sc_hd__and4_1 _10708_ (.A(_04837_),
    .B(_04843_),
    .C(_04857_),
    .D(_04869_),
    .X(_04874_));
 sky130_fd_sc_hd__nor2_1 _10709_ (.A(_04862_),
    .B(_04869_),
    .Y(_04875_));
 sky130_fd_sc_hd__o31a_1 _10710_ (.A1(_04874_),
    .A2(_04875_),
    .A3(net100),
    .B1(_04643_),
    .X(_04876_));
 sky130_fd_sc_hd__a22oi_1 _10711_ (.A1(_04873_),
    .A2(_04876_),
    .B1(_04867_),
    .B2(_03603_),
    .Y(net88));
 sky130_fd_sc_hd__a41o_1 _10712_ (.A1(_04583_),
    .A2(_04830_),
    .A3(_04858_),
    .A4(_04870_),
    .B1(_03610_),
    .X(_04878_));
 sky130_fd_sc_hd__a41oi_1 _10713_ (.A1(_04832_),
    .A2(_04870_),
    .A3(_04858_),
    .A4(_03610_),
    .B1(_04572_),
    .Y(_04879_));
 sky130_fd_sc_hd__and3_1 _10714_ (.A(_03610_),
    .B(_04862_),
    .C(_04869_),
    .X(_04880_));
 sky130_fd_sc_hd__o2bb2a_1 _10715_ (.A1_N(_04862_),
    .A2_N(_04869_),
    .B1(net24),
    .B2(net56),
    .X(_04881_));
 sky130_fd_sc_hd__o31ai_1 _10716_ (.A1(_04880_),
    .A2(_04881_),
    .A3(net100),
    .B1(_04636_),
    .Y(_04882_));
 sky130_fd_sc_hd__a21oi_1 _10717_ (.A1(_04879_),
    .A2(_04878_),
    .B1(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__a41oi_1 _10718_ (.A1(_01375_),
    .A2(_01507_),
    .A3(_03556_),
    .A4(_03565_),
    .B1(_03587_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand4_1 _10719_ (.A(_03556_),
    .B(_03565_),
    .C(_03571_),
    .D(_03587_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_1 _10720_ (.A1(_01518_),
    .A2(_04885_),
    .B1(_03612_),
    .Y(_04886_));
 sky130_fd_sc_hd__o21ai_1 _10721_ (.A1(_04884_),
    .A2(_04886_),
    .B1(_03598_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand2_1 _10722_ (.A(_04888_),
    .B(_03600_),
    .Y(_04889_));
 sky130_fd_sc_hd__a2bb2oi_1 _10723_ (.A1_N(_04644_),
    .A2_N(_04883_),
    .B1(_04889_),
    .B2(_03603_),
    .Y(net90));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(net57),
    .A1(net25),
    .S(net102),
    .X(_04890_));
 sky130_fd_sc_hd__nand3_1 _10725_ (.A(_04636_),
    .B(_04890_),
    .C(_03601_),
    .Y(_04891_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(net25),
    .A1(net57),
    .S(_00803_),
    .X(_04892_));
 sky130_fd_sc_hd__nand2_1 _10727_ (.A(_03602_),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__o311a_1 _10728_ (.A1(_00803_),
    .A2(_00891_),
    .A3(_03618_),
    .B1(_00748_),
    .C1(_05339_),
    .X(_04894_));
 sky130_fd_sc_hd__a21bo_1 _10729_ (.A1(_04891_),
    .A2(_04893_),
    .B1_N(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__o31ai_1 _10730_ (.A1(_00935_),
    .A2(_03599_),
    .A3(_03618_),
    .B1(_04895_),
    .Y(net91));
 sky130_fd_sc_hd__a41o_1 _10731_ (.A1(_03592_),
    .A2(_03594_),
    .A3(_03572_),
    .A4(_03573_),
    .B1(_05339_),
    .X(_04897_));
 sky130_fd_sc_hd__o21a_1 _10732_ (.A1(net65),
    .A2(_04572_),
    .B1(_04897_),
    .X(net66));
 sky130_fd_sc_hd__buf_12 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_16 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_16 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_16 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_16 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_16 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_12 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_12 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_12 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_12 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_16 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_12 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_12 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_16 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_12 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_12 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_12 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_16 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_16 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_16 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_16 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_16 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_6 input65 (.A(sel),
    .X(net65));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(overflow));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(result[0]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(result[10]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(result[11]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(result[12]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(result[13]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(result[14]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(result[15]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(result[16]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(result[17]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(result[18]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(result[19]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(result[1]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(result[20]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(result[21]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(result[22]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(result[23]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(result[24]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(result[25]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(result[26]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(result[27]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(result[28]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(result[29]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(result[2]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(result[30]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(result[31]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(result[3]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(result[4]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(result[5]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(result[6]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(result[7]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(result[8]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(result[9]));
 sky130_fd_sc_hd__buf_12 max_cap99 (.A(_03606_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_8 max_cap100 (.A(_04573_),
    .X(net100));
 sky130_fd_sc_hd__buf_12 max_cap101 (.A(_04256_),
    .X(net101));
 sky130_fd_sc_hd__buf_12 max_cap102 (.A(_04256_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 max_cap103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_4 max_cap104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 max_cap105 (.A(_03611_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_16 max_cap106 (.A(_03731_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_8 max_cap107 (.A(_03737_),
    .X(net107));
 sky130_fd_sc_hd__buf_12 max_cap108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_8 max_cap109 (.A(_03651_),
    .X(net109));
 sky130_fd_sc_hd__buf_12 max_cap110 (.A(_03642_),
    .X(net110));
 sky130_fd_sc_hd__buf_12 max_cap111 (.A(_03642_),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 max_cap112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 max_cap113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__buf_4 max_cap114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_8 max_cap115 (.A(_03650_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_16 max_cap116 (.A(_00880_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_16 wire117 (.A(_00792_),
    .X(net117));
 sky130_fd_sc_hd__buf_4 wire118 (.A(_00836_),
    .X(net118));
endmodule
